// carry_lookahead_toplayici.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module carry_lookahead_toplayici(


);


endmodule
