
`include "tanimlamalar.vh"

`ifndef OPENLANE
module toplayici(
	input  [32:0] a_in,
	input  [32:0] b_in,
	output [32:0] sum
);
	wire n8_tree_32, n9_tree_32, n10_tree_32, n11_tree_32, n12_tree_32, n13_tree_32, n16_tree_32, n17_tree_32, n18_tree_31, n18_tree_32, n19_tree_31, n19_tree_32, n20_tree_32, n21_tree_32, n24_tree_32, n25_tree_32, n26_tree_32, n27_tree_32, n28_tree_32, n29_tree_32, n32_tree_32, n33_tree_32, n34_tree_31, n34_tree_32, n35_tree_31, n35_tree_32, n36_tree_32, n37_tree_32, n38_tree_30, n39_tree_30, n40_tree_32, n41_tree_32, n42_tree_32, n43_tree_32, n44_tree_32, n45_tree_32, n48_tree_32, n49_tree_32, n50_tree_31, n50_tree_32, n51_tree_31, n51_tree_32, n52_tree_32, n53_tree_32, n56_tree_32, n57_tree_32, n58_tree_32, n59_tree_32, n60_tree_32, n61_tree_32, n64_tree_32, n65_tree_32, n66_tree_31, n66_tree_32, n67_tree_31, n67_tree_32, n68_tree_32, n69_tree_32, n70_tree_30, n71_tree_30, n72_tree_32, n73_tree_32, n74_tree_32, n75_tree_32, n76_tree_32, n77_tree_32, n80_tree_32, n81_tree_32, n82_tree_31, n82_tree_32, n83_tree_31, n83_tree_32, n84_tree_32, n85_tree_32, n88_tree_32, n89_tree_32, n90_tree_32, n91_tree_32, n92_tree_32, n93_tree_32, n96_tree_32, n97_tree_32, n98_tree_31, n98_tree_32, n99_tree_31, n99_tree_32, n100_tree_32, n101_tree_32, n104_tree_32, n105_tree_32, n106_tree_32, n107_tree_32, n108_tree_32, n109_tree_32, n112_tree_32, n113_tree_32, n114_tree_28, n114_tree_32, n115_tree_32, n116_tree_32, n117_tree_32, n119_tree_29, n120_tree_32, n121_tree_32, n124_tree_30, n124_tree_32, n125_tree_32, n129_tree_31, n134_tree_32;

	adder_tree_32 U0(
		.a_in(a_in[32:0]),
		.b_in(b_in[32:0]),
		.sum(sum[32]),
		.n125_tree_32(n125_tree_32),
		.n124_tree_32(n124_tree_32),
		.n121_tree_32(n121_tree_32),
		.n120_tree_32(n120_tree_32),
		.n117_tree_32(n117_tree_32),
		.n116_tree_32(n116_tree_32),
		.n113_tree_32(n113_tree_32),
		.n112_tree_32(n112_tree_32),
		.n109_tree_32(n109_tree_32),
		.n108_tree_32(n108_tree_32),
		.n105_tree_32(n105_tree_32),
		.n104_tree_32(n104_tree_32),
		.n101_tree_32(n101_tree_32),
		.n100_tree_32(n100_tree_32),
		.n97_tree_32(n97_tree_32),
		.n96_tree_32(n96_tree_32),
		.n93_tree_32(n93_tree_32),
		.n92_tree_32(n92_tree_32),
		.n89_tree_32(n89_tree_32),
		.n88_tree_32(n88_tree_32),
		.n85_tree_32(n85_tree_32),
		.n84_tree_32(n84_tree_32),
		.n81_tree_32(n81_tree_32),
		.n80_tree_32(n80_tree_32),
		.n77_tree_32(n77_tree_32),
		.n76_tree_32(n76_tree_32),
		.n73_tree_32(n73_tree_32),
		.n72_tree_32(n72_tree_32),
		.n69_tree_32(n69_tree_32),
		.n68_tree_32(n68_tree_32),
		.n65_tree_32(n65_tree_32),
		.n64_tree_32(n64_tree_32),
		.n61_tree_32(n61_tree_32),
		.n60_tree_32(n60_tree_32),
		.n57_tree_32(n57_tree_32),
		.n56_tree_32(n56_tree_32),
		.n53_tree_32(n53_tree_32),
		.n52_tree_32(n52_tree_32),
		.n49_tree_32(n49_tree_32),
		.n48_tree_32(n48_tree_32),
		.n45_tree_32(n45_tree_32),
		.n44_tree_32(n44_tree_32),
		.n41_tree_32(n41_tree_32),
		.n40_tree_32(n40_tree_32),
		.n37_tree_32(n37_tree_32),
		.n36_tree_32(n36_tree_32),
		.n33_tree_32(n33_tree_32),
		.n32_tree_32(n32_tree_32),
		.n29_tree_32(n29_tree_32),
		.n28_tree_32(n28_tree_32),
		.n25_tree_32(n25_tree_32),
		.n24_tree_32(n24_tree_32),
		.n21_tree_32(n21_tree_32),
		.n20_tree_32(n20_tree_32),
		.n17_tree_32(n17_tree_32),
		.n16_tree_32(n16_tree_32),
		.n13_tree_32(n13_tree_32),
		.n12_tree_32(n12_tree_32),
		.n9_tree_32(n9_tree_32),
		.n8_tree_32(n8_tree_32),
		.n10_tree_32(n10_tree_32),
		.n11_tree_32(n11_tree_32),
		.n18_tree_32(n18_tree_32),
		.n19_tree_32(n19_tree_32),
		.n26_tree_32(n26_tree_32),
		.n27_tree_32(n27_tree_32),
		.n34_tree_32(n34_tree_32),
		.n35_tree_32(n35_tree_32),
		.n42_tree_32(n42_tree_32),
		.n43_tree_32(n43_tree_32),
		.n50_tree_32(n50_tree_32),
		.n51_tree_32(n51_tree_32),
		.n58_tree_32(n58_tree_32),
		.n59_tree_32(n59_tree_32),
		.n66_tree_32(n66_tree_32),
		.n67_tree_32(n67_tree_32),
		.n74_tree_32(n74_tree_32),
		.n75_tree_32(n75_tree_32),
		.n82_tree_32(n82_tree_32),
		.n83_tree_32(n83_tree_32),
		.n90_tree_32(n90_tree_32),
		.n91_tree_32(n91_tree_32),
		.n98_tree_32(n98_tree_32),
		.n99_tree_32(n99_tree_32),
		.n106_tree_32(n106_tree_32),
		.n107_tree_32(n107_tree_32),
		.n114_tree_32(n114_tree_32),
		.n115_tree_32(n115_tree_32),
		.n134_tree_32(n134_tree_32)
	);
	adder_tree_31 U1(
		.a_in(a_in[31:0]),
		.b_in(b_in[31:0]),
		.n125_tree_32(n125_tree_32),
		.n124_tree_32(n124_tree_32),
		.n9_tree_32(n9_tree_32),
		.n8_tree_32(n8_tree_32),
		.n10_tree_32(n10_tree_32),
		.n11_tree_32(n11_tree_32),
		.n18_tree_32(n18_tree_32),
		.n19_tree_32(n19_tree_32),
		.n26_tree_32(n26_tree_32),
		.n27_tree_32(n27_tree_32),
		.n34_tree_32(n34_tree_32),
		.n35_tree_32(n35_tree_32),
		.n42_tree_32(n42_tree_32),
		.n43_tree_32(n43_tree_32),
		.n50_tree_32(n50_tree_32),
		.n51_tree_32(n51_tree_32),
		.n58_tree_32(n58_tree_32),
		.n59_tree_32(n59_tree_32),
		.n66_tree_32(n66_tree_32),
		.n67_tree_32(n67_tree_32),
		.n74_tree_32(n74_tree_32),
		.n75_tree_32(n75_tree_32),
		.n82_tree_32(n82_tree_32),
		.n83_tree_32(n83_tree_32),
		.n90_tree_32(n90_tree_32),
		.n91_tree_32(n91_tree_32),
		.n98_tree_32(n98_tree_32),
		.n99_tree_32(n99_tree_32),
		.n106_tree_32(n106_tree_32),
		.n107_tree_32(n107_tree_32),
		.n114_tree_32(n114_tree_32),
		.n115_tree_32(n115_tree_32),
		.n134_tree_32(n134_tree_32),
		.sum(sum[31]),
		.n18_tree_31(n18_tree_31),
		.n19_tree_31(n19_tree_31),
		.n34_tree_31(n34_tree_31),
		.n35_tree_31(n35_tree_31),
		.n50_tree_31(n50_tree_31),
		.n51_tree_31(n51_tree_31),
		.n66_tree_31(n66_tree_31),
		.n67_tree_31(n67_tree_31),
		.n82_tree_31(n82_tree_31),
		.n83_tree_31(n83_tree_31),
		.n98_tree_31(n98_tree_31),
		.n99_tree_31(n99_tree_31),
		.n129_tree_31(n129_tree_31)
	);
	adder_tree_30 U2(
		.a_in(a_in[30:0]),
		.b_in(b_in[30:0]),
		.n10_tree_32(n10_tree_32),
		.n11_tree_32(n11_tree_32),
		.n18_tree_31(n18_tree_31),
		.n19_tree_31(n19_tree_31),
		.n34_tree_31(n34_tree_31),
		.n35_tree_31(n35_tree_31),
		.n50_tree_31(n50_tree_31),
		.n51_tree_31(n51_tree_31),
		.n66_tree_31(n66_tree_31),
		.n67_tree_31(n67_tree_31),
		.n82_tree_31(n82_tree_31),
		.n83_tree_31(n83_tree_31),
		.n98_tree_31(n98_tree_31),
		.n99_tree_31(n99_tree_31),
		.n114_tree_32(n114_tree_32),
		.n115_tree_32(n115_tree_32),
		.n129_tree_31(n129_tree_31),
		.sum(sum[30]),
		.n38_tree_30(n38_tree_30),
		.n39_tree_30(n39_tree_30),
		.n70_tree_30(n70_tree_30),
		.n71_tree_30(n71_tree_30),
		.n124_tree_30(n124_tree_30)
	);
	adder_tree_29 U3(
		.a_in(a_in[29:0]),
		.b_in(b_in[29:0]),
		.n17_tree_32(n17_tree_32),
		.n16_tree_32(n16_tree_32),
		.n18_tree_31(n18_tree_31),
		.n19_tree_31(n19_tree_31),
		.n38_tree_30(n38_tree_30),
		.n39_tree_30(n39_tree_30),
		.n70_tree_30(n70_tree_30),
		.n71_tree_30(n71_tree_30),
		.n98_tree_31(n98_tree_31),
		.n99_tree_31(n99_tree_31),
		.n124_tree_30(n124_tree_30),
		.sum(sum[29]),
		.n119_tree_29(n119_tree_29)
	);
	adder_tree_28 U4(
		.a_in(a_in[28:0]),
		.b_in(b_in[28:0]),
		.n18_tree_31(n18_tree_31),
		.n19_tree_31(n19_tree_31),
		.n38_tree_30(n38_tree_30),
		.n39_tree_30(n39_tree_30),
		.n70_tree_30(n70_tree_30),
		.n71_tree_30(n71_tree_30),
		.n119_tree_29(n119_tree_29),
		.sum(sum[28]),
		.n114_tree_28(n114_tree_28)
	);
	adder_tree_27 U5(
		.a_in(a_in[27:0]),
		.b_in(b_in[27:0]),
		.n25_tree_32(n25_tree_32),
		.n24_tree_32(n24_tree_32),
		.n26_tree_32(n26_tree_32),
		.n27_tree_32(n27_tree_32),
		.n38_tree_30(n38_tree_30),
		.n39_tree_30(n39_tree_30),
		.n114_tree_28(n114_tree_28),
		.sum(sum[27])
	);
	adder_tree_26 U6(
		.a_in(a_in[26:0]),
		.b_in(b_in[26:0]),
		.n26_tree_32(n26_tree_32),
		.n27_tree_32(n27_tree_32),
		.n38_tree_30(n38_tree_30),
		.n39_tree_30(n39_tree_30),
		.n114_tree_28(n114_tree_28),
		.sum(sum[26])
	);
	adder_tree_25 U7(
		.a_in(a_in[25:0]),
		.b_in(b_in[25:0]),
		.n33_tree_32(n33_tree_32),
		.n32_tree_32(n32_tree_32),
		.n38_tree_30(n38_tree_30),
		.n39_tree_30(n39_tree_30),
		.n114_tree_28(n114_tree_28),
		.sum(sum[25])
	);
	adder_tree_24 U8(
		.a_in(a_in[24:0]),
		.b_in(b_in[24:0]),
		.n38_tree_30(n38_tree_30),
		.n39_tree_30(n39_tree_30),
		.n114_tree_28(n114_tree_28),
		.sum(sum[24])
	);
	adder_tree_23 U9(
		.a_in(a_in[23:0]),
		.b_in(b_in[23:0]),
		.n41_tree_32(n41_tree_32),
		.n40_tree_32(n40_tree_32),
		.n42_tree_32(n42_tree_32),
		.n43_tree_32(n43_tree_32),
		.n50_tree_31(n50_tree_31),
		.n51_tree_31(n51_tree_31),
		.n114_tree_28(n114_tree_28),
		.sum(sum[23])
	);
	adder_tree_22 U10(
		.a_in(a_in[22:0]),
		.b_in(b_in[22:0]),
		.n42_tree_32(n42_tree_32),
		.n43_tree_32(n43_tree_32),
		.n50_tree_31(n50_tree_31),
		.n51_tree_31(n51_tree_31),
		.n114_tree_28(n114_tree_28),
		.sum(sum[22])
	);
	adder_tree_21 U11(
		.a_in(a_in[21:0]),
		.b_in(b_in[21:0]),
		.n49_tree_32(n49_tree_32),
		.n48_tree_32(n48_tree_32),
		.n50_tree_31(n50_tree_31),
		.n51_tree_31(n51_tree_31),
		.n114_tree_28(n114_tree_28),
		.sum(sum[21])
	);
	adder_tree_20 U12(
		.a_in(a_in[20:0]),
		.b_in(b_in[20:0]),
		.n50_tree_31(n50_tree_31),
		.n51_tree_31(n51_tree_31),
		.n114_tree_28(n114_tree_28),
		.sum(sum[20])
	);
	adder_tree_19 U13(
		.a_in(a_in[19:0]),
		.b_in(b_in[19:0]),
		.n57_tree_32(n57_tree_32),
		.n56_tree_32(n56_tree_32),
		.n58_tree_32(n58_tree_32),
		.n59_tree_32(n59_tree_32),
		.n114_tree_28(n114_tree_28),
		.sum(sum[19])
	);
	adder_tree_18 U14(
		.a_in(a_in[18:0]),
		.b_in(b_in[18:0]),
		.n58_tree_32(n58_tree_32),
		.n59_tree_32(n59_tree_32),
		.n114_tree_28(n114_tree_28),
		.sum(sum[18])
	);
	adder_tree_17 U15(
		.a_in(a_in[17:0]),
		.b_in(b_in[17:0]),
		.n65_tree_32(n65_tree_32),
		.n64_tree_32(n64_tree_32),
		.n114_tree_28(n114_tree_28),
		.sum(sum[17])
	);
	adder_tree_16 U16(
		.a_in(a_in[16:0]),
		.b_in(b_in[16:0]),
		.n114_tree_28(n114_tree_28),
		.sum(sum[16])
	);
	adder_tree_15 U17(
		.a_in(a_in[15:0]),
		.b_in(b_in[15:0]),
		.n73_tree_32(n73_tree_32),
		.n72_tree_32(n72_tree_32),
		.n74_tree_32(n74_tree_32),
		.n75_tree_32(n75_tree_32),
		.n82_tree_31(n82_tree_31),
		.n83_tree_31(n83_tree_31),
		.n119_tree_29(n119_tree_29),
		.sum(sum[15])
	);
	adder_tree_14 U18(
		.a_in(a_in[14:0]),
		.b_in(b_in[14:0]),
		.n74_tree_32(n74_tree_32),
		.n75_tree_32(n75_tree_32),
		.n82_tree_31(n82_tree_31),
		.n83_tree_31(n83_tree_31),
		.n119_tree_29(n119_tree_29),
		.sum(sum[14])
	);
	adder_tree_13 U19(
		.a_in(a_in[13:0]),
		.b_in(b_in[13:0]),
		.n81_tree_32(n81_tree_32),
		.n80_tree_32(n80_tree_32),
		.n82_tree_31(n82_tree_31),
		.n83_tree_31(n83_tree_31),
		.n119_tree_29(n119_tree_29),
		.sum(sum[13])
	);
	adder_tree_12 U20(
		.a_in(a_in[12:0]),
		.b_in(b_in[12:0]),
		.n82_tree_31(n82_tree_31),
		.n83_tree_31(n83_tree_31),
		.n119_tree_29(n119_tree_29),
		.sum(sum[12])
	);
	adder_tree_11 U21(
		.a_in(a_in[11:0]),
		.b_in(b_in[11:0]),
		.n89_tree_32(n89_tree_32),
		.n88_tree_32(n88_tree_32),
		.n90_tree_32(n90_tree_32),
		.n91_tree_32(n91_tree_32),
		.n119_tree_29(n119_tree_29),
		.sum(sum[11])
	);
	adder_tree_10 U22(
		.a_in(a_in[10:0]),
		.b_in(b_in[10:0]),
		.n90_tree_32(n90_tree_32),
		.n91_tree_32(n91_tree_32),
		.n119_tree_29(n119_tree_29),
		.sum(sum[10])
	);
	adder_tree_9 U23(
		.a_in(a_in[9:0]),
		.b_in(b_in[9:0]),
		.n97_tree_32(n97_tree_32),
		.n96_tree_32(n96_tree_32),
		.n119_tree_29(n119_tree_29),
		.sum(sum[9])
	);
	adder_tree_8 U24(
		.a_in(a_in[8:0]),
		.b_in(b_in[8:0]),
		.n119_tree_29(n119_tree_29),
		.sum(sum[8])
	);
	adder_tree_7 U25(
		.a_in(a_in[7:0]),
		.b_in(b_in[7:0]),
		.n105_tree_32(n105_tree_32),
		.n104_tree_32(n104_tree_32),
		.n106_tree_32(n106_tree_32),
		.n107_tree_32(n107_tree_32),
		.n124_tree_30(n124_tree_30),
		.sum(sum[7])
	);
	adder_tree_6 U26(
		.a_in(a_in[6:0]),
		.b_in(b_in[6:0]),
		.n106_tree_32(n106_tree_32),
		.n107_tree_32(n107_tree_32),
		.n124_tree_30(n124_tree_30),
		.sum(sum[6])
	);
	adder_tree_5 U27(
		.a_in(a_in[5:0]),
		.b_in(b_in[5:0]),
		.n113_tree_32(n113_tree_32),
		.n112_tree_32(n112_tree_32),
		.n124_tree_30(n124_tree_30),
		.sum(sum[5])
	);
	adder_tree_4 U28(
		.a_in(a_in[4:0]),
		.b_in(b_in[4:0]),
		.n124_tree_30(n124_tree_30),
		.sum(sum[4])
	);
	adder_tree_3 U29(
		.a_in(a_in[3:0]),
		.b_in(b_in[3:0]),
		.n121_tree_32(n121_tree_32),
		.n120_tree_32(n120_tree_32),
		.n129_tree_31(n129_tree_31),
		.sum(sum[3])
	);
	adder_tree_2 U30(
		.a_in(a_in[2:0]),
		.b_in(b_in[2:0]),
		.n129_tree_31(n129_tree_31),
		.sum(sum[2])
	);
	adder_tree_1 U31(
		.a_in(a_in[1:0]),
		.b_in(b_in[1:0]),
		.n134_tree_32(n134_tree_32),
		.sum(sum[1])
	);
	adder_tree_0 U32(
		.a_in(a_in[0]),
		.b_in(b_in[0]),
		.sum(sum[0])
	);
endmodule // adder
module adder_tree_0(
	input   a_in,
	input   b_in,
	output  sum
);
// adder_forest tree_0
	wire n1_tree_0;
	assign sum = n1_tree_0;
    assign n1_tree_0 = a_in^b_in;
endmodule // adder_tree_0
module adder_tree_1(
	input  [1:0] a_in,
	input  [1:0] b_in,
	input   n134_tree_32,
	output  sum
);
// adder_forest tree_1
	wire n5_tree_1;
    assign sum = n134_tree_32^n5_tree_1;
    assign n5_tree_1 = a_in[1]^b_in[1];
endmodule // adder_tree_1
module adder_tree_2(
	input  [2:0] a_in,
	input  [2:0] b_in,
	input   n129_tree_31,
	output  sum
);
// adder_forest tree_2
	wire n10_tree_2;
    assign sum = n129_tree_31^n10_tree_2;
    assign n10_tree_2 = a_in[2]^b_in[2];
endmodule // adder_tree_2
module adder_tree_3(
	input  [3:0] a_in,
	input  [3:0] b_in,
	input   n121_tree_32,
	input   n120_tree_32,
	input   n129_tree_31,
	output  sum
);
// adder_forest tree_3
	wire n12_tree_3, n15_tree_3;
    assign n12_tree_3 = (n129_tree_31&n121_tree_32)|n120_tree_32;
    assign sum = n12_tree_3^n15_tree_3;
    assign n15_tree_3 = a_in[3]^b_in[3];
endmodule // adder_tree_3
module adder_tree_4(
	input  [4:0] a_in,
	input  [4:0] b_in,
	input   n124_tree_30,
	output  sum
);
// adder_forest tree_4
	wire n20_tree_4;
    assign sum = n124_tree_30^n20_tree_4;
    assign n20_tree_4 = a_in[4]^b_in[4];
endmodule // adder_tree_4
module adder_tree_5(
	input  [5:0] a_in,
	input  [5:0] b_in,
	input   n113_tree_32,
	input   n112_tree_32,
	input   n124_tree_30,
	output  sum
);
// adder_forest tree_5
	wire n20_tree_5, n24_tree_5;
    assign n20_tree_5 = (n124_tree_30&n113_tree_32)|n112_tree_32;
    assign sum = n20_tree_5^n24_tree_5;
    assign n24_tree_5 = a_in[5]^b_in[5];
endmodule // adder_tree_5
module adder_tree_6(
	input  [6:0] a_in,
	input  [6:0] b_in,
	input   n106_tree_32,
	input   n107_tree_32,
	input   n124_tree_30,
	output  sum
);
// adder_forest tree_6
	wire n25_tree_6, n29_tree_6;
    assign n25_tree_6 = (n124_tree_30&n107_tree_32)|n106_tree_32;
    assign sum = n25_tree_6^n29_tree_6;
    assign n29_tree_6 = a_in[6]^b_in[6];
endmodule // adder_tree_6
module adder_tree_7(
	input  [7:0] a_in,
	input  [7:0] b_in,
	input   n105_tree_32,
	input   n104_tree_32,
	input   n106_tree_32,
	input   n107_tree_32,
	input   n124_tree_30,
	output  sum
);
// adder_forest tree_7
	wire n3_tree_7, n28_tree_7, n29_tree_7, n33_tree_7;
    assign n28_tree_7 = n105_tree_32&n107_tree_32;
    assign n3_tree_7 = (n106_tree_32&n105_tree_32)|n104_tree_32;
    assign n29_tree_7 = (n124_tree_30&n28_tree_7)|n3_tree_7;
    assign sum = n29_tree_7^n33_tree_7;
    assign n33_tree_7 = a_in[7]^b_in[7];
endmodule // adder_tree_7
module adder_tree_8(
	input  [8:0] a_in,
	input  [8:0] b_in,
	input   n119_tree_29,
	output  sum
);
// adder_forest tree_8
	wire n37_tree_8;
    assign sum = n119_tree_29^n37_tree_8;
    assign n37_tree_8 = a_in[8]^b_in[8];
endmodule // adder_tree_8
module adder_tree_9(
	input  [9:0] a_in,
	input  [9:0] b_in,
	input   n97_tree_32,
	input   n96_tree_32,
	input   n119_tree_29,
	output  sum
);
// adder_forest tree_9
	wire n36_tree_9, n41_tree_9;
    assign n36_tree_9 = (n119_tree_29&n97_tree_32)|n96_tree_32;
    assign sum = n36_tree_9^n41_tree_9;
    assign n41_tree_9 = a_in[9]^b_in[9];
endmodule // adder_tree_9
module adder_tree_10(
	input  [10:0] a_in,
	input  [10:0] b_in,
	input   n90_tree_32,
	input   n91_tree_32,
	input   n119_tree_29,
	output  sum
);
// adder_forest tree_10
	wire n41_tree_10, n46_tree_10;
    assign n41_tree_10 = (n119_tree_29&n91_tree_32)|n90_tree_32;
    assign sum = n41_tree_10^n46_tree_10;
    assign n46_tree_10 = a_in[10]^b_in[10];
endmodule // adder_tree_10
module adder_tree_11(
	input  [11:0] a_in,
	input  [11:0] b_in,
	input   n89_tree_32,
	input   n88_tree_32,
	input   n90_tree_32,
	input   n91_tree_32,
	input   n119_tree_29,
	output  sum
);
// adder_forest tree_11
	wire n3_tree_11, n44_tree_11, n45_tree_11, n50_tree_11;
    assign n44_tree_11 = n89_tree_32&n91_tree_32;
    assign n3_tree_11 = (n90_tree_32&n89_tree_32)|n88_tree_32;
    assign n45_tree_11 = (n119_tree_29&n44_tree_11)|n3_tree_11;
    assign sum = n45_tree_11^n50_tree_11;
    assign n50_tree_11 = a_in[11]^b_in[11];
endmodule // adder_tree_11
module adder_tree_12(
	input  [12:0] a_in,
	input  [12:0] b_in,
	input   n82_tree_31,
	input   n83_tree_31,
	input   n119_tree_29,
	output  sum
);
// adder_forest tree_12
	wire n49_tree_12, n54_tree_12;
    assign n49_tree_12 = (n119_tree_29&n83_tree_31)|n82_tree_31;
    assign sum = n49_tree_12^n54_tree_12;
    assign n54_tree_12 = a_in[12]^b_in[12];
endmodule // adder_tree_12
module adder_tree_13(
	input  [13:0] a_in,
	input  [13:0] b_in,
	input   n81_tree_32,
	input   n80_tree_32,
	input   n82_tree_31,
	input   n83_tree_31,
	input   n119_tree_29,
	output  sum
);
// adder_forest tree_13
	wire n3_tree_13, n52_tree_13, n53_tree_13, n58_tree_13;
    assign n52_tree_13 = n81_tree_32&n83_tree_31;
    assign n3_tree_13 = (n82_tree_31&n81_tree_32)|n80_tree_32;
    assign n53_tree_13 = (n119_tree_29&n52_tree_13)|n3_tree_13;
    assign sum = n53_tree_13^n58_tree_13;
    assign n58_tree_13 = a_in[13]^b_in[13];
endmodule // adder_tree_13
module adder_tree_14(
	input  [14:0] a_in,
	input  [14:0] b_in,
	input   n74_tree_32,
	input   n75_tree_32,
	input   n82_tree_31,
	input   n83_tree_31,
	input   n119_tree_29,
	output  sum
);
// adder_forest tree_14
	wire n6_tree_14, n7_tree_14, n57_tree_14, n62_tree_14;
    assign n7_tree_14 = n75_tree_32&n83_tree_31;
    assign n6_tree_14 = (n82_tree_31&n75_tree_32)|n74_tree_32;
    assign n57_tree_14 = (n119_tree_29&n7_tree_14)|n6_tree_14;
    assign sum = n57_tree_14^n62_tree_14;
    assign n62_tree_14 = a_in[14]^b_in[14];
endmodule // adder_tree_14
module adder_tree_15(
	input  [15:0] a_in,
	input  [15:0] b_in,
	input   n73_tree_32,
	input   n72_tree_32,
	input   n74_tree_32,
	input   n75_tree_32,
	input   n82_tree_31,
	input   n83_tree_31,
	input   n119_tree_29,
	output  sum
);
// adder_forest tree_15
	wire n3_tree_15, n10_tree_15, n11_tree_15, n60_tree_15, n61_tree_15, n66_tree_15;
    assign n60_tree_15 = n73_tree_32&n75_tree_32;
    assign n3_tree_15 = (n74_tree_32&n73_tree_32)|n72_tree_32;
    assign n11_tree_15 = n60_tree_15&n83_tree_31;
    assign n10_tree_15 = (n82_tree_31&n60_tree_15)|n3_tree_15;
    assign n61_tree_15 = (n119_tree_29&n11_tree_15)|n10_tree_15;
    assign sum = n61_tree_15^n66_tree_15;
    assign n66_tree_15 = a_in[15]^b_in[15];
endmodule // adder_tree_15
module adder_tree_16(
	input  [16:0] a_in,
	input  [16:0] b_in,
	input   n114_tree_28,
	output  sum
);
// adder_forest tree_16
	wire n70_tree_16;
    assign sum = n114_tree_28^n70_tree_16;
    assign n70_tree_16 = a_in[16]^b_in[16];
endmodule // adder_tree_16
module adder_tree_17(
	input  [17:0] a_in,
	input  [17:0] b_in,
	input   n65_tree_32,
	input   n64_tree_32,
	input   n114_tree_28,
	output  sum
);
// adder_forest tree_17
	wire n68_tree_17, n74_tree_17;
    assign n68_tree_17 = (n114_tree_28&n65_tree_32)|n64_tree_32;
    assign sum = n68_tree_17^n74_tree_17;
    assign n74_tree_17 = a_in[17]^b_in[17];
endmodule // adder_tree_17
module adder_tree_18(
	input  [18:0] a_in,
	input  [18:0] b_in,
	input   n58_tree_32,
	input   n59_tree_32,
	input   n114_tree_28,
	output  sum
);
// adder_forest tree_18
	wire n73_tree_18, n79_tree_18;
    assign n73_tree_18 = (n114_tree_28&n59_tree_32)|n58_tree_32;
    assign sum = n73_tree_18^n79_tree_18;
    assign n79_tree_18 = a_in[18]^b_in[18];
endmodule // adder_tree_18
module adder_tree_19(
	input  [19:0] a_in,
	input  [19:0] b_in,
	input   n57_tree_32,
	input   n56_tree_32,
	input   n58_tree_32,
	input   n59_tree_32,
	input   n114_tree_28,
	output  sum
);
// adder_forest tree_19
	wire n3_tree_19, n76_tree_19, n77_tree_19, n83_tree_19;
    assign n76_tree_19 = n57_tree_32&n59_tree_32;
    assign n3_tree_19 = (n58_tree_32&n57_tree_32)|n56_tree_32;
    assign n77_tree_19 = (n114_tree_28&n76_tree_19)|n3_tree_19;
    assign sum = n77_tree_19^n83_tree_19;
    assign n83_tree_19 = a_in[19]^b_in[19];
endmodule // adder_tree_19
module adder_tree_20(
	input  [20:0] a_in,
	input  [20:0] b_in,
	input   n50_tree_31,
	input   n51_tree_31,
	input   n114_tree_28,
	output  sum
);
// adder_forest tree_20
	wire n81_tree_20, n87_tree_20;
    assign n81_tree_20 = (n114_tree_28&n51_tree_31)|n50_tree_31;
    assign sum = n81_tree_20^n87_tree_20;
    assign n87_tree_20 = a_in[20]^b_in[20];
endmodule // adder_tree_20
module adder_tree_21(
	input  [21:0] a_in,
	input  [21:0] b_in,
	input   n49_tree_32,
	input   n48_tree_32,
	input   n50_tree_31,
	input   n51_tree_31,
	input   n114_tree_28,
	output  sum
);
// adder_forest tree_21
	wire n3_tree_21, n84_tree_21, n85_tree_21, n91_tree_21;
    assign n84_tree_21 = n49_tree_32&n51_tree_31;
    assign n3_tree_21 = (n50_tree_31&n49_tree_32)|n48_tree_32;
    assign n85_tree_21 = (n114_tree_28&n84_tree_21)|n3_tree_21;
    assign sum = n85_tree_21^n91_tree_21;
    assign n91_tree_21 = a_in[21]^b_in[21];
endmodule // adder_tree_21
module adder_tree_22(
	input  [22:0] a_in,
	input  [22:0] b_in,
	input   n42_tree_32,
	input   n43_tree_32,
	input   n50_tree_31,
	input   n51_tree_31,
	input   n114_tree_28,
	output  sum
);
// adder_forest tree_22
	wire n6_tree_22, n7_tree_22, n89_tree_22, n95_tree_22;
    assign n7_tree_22 = n43_tree_32&n51_tree_31;
    assign n6_tree_22 = (n50_tree_31&n43_tree_32)|n42_tree_32;
    assign n89_tree_22 = (n114_tree_28&n7_tree_22)|n6_tree_22;
    assign sum = n89_tree_22^n95_tree_22;
    assign n95_tree_22 = a_in[22]^b_in[22];
endmodule // adder_tree_22
module adder_tree_23(
	input  [23:0] a_in,
	input  [23:0] b_in,
	input   n41_tree_32,
	input   n40_tree_32,
	input   n42_tree_32,
	input   n43_tree_32,
	input   n50_tree_31,
	input   n51_tree_31,
	input   n114_tree_28,
	output  sum
);
// adder_forest tree_23
	wire n3_tree_23, n10_tree_23, n11_tree_23, n92_tree_23, n93_tree_23, n99_tree_23;
    assign n92_tree_23 = n41_tree_32&n43_tree_32;
    assign n3_tree_23 = (n42_tree_32&n41_tree_32)|n40_tree_32;
    assign n11_tree_23 = n92_tree_23&n51_tree_31;
    assign n10_tree_23 = (n50_tree_31&n92_tree_23)|n3_tree_23;
    assign n93_tree_23 = (n114_tree_28&n11_tree_23)|n10_tree_23;
    assign sum = n93_tree_23^n99_tree_23;
    assign n99_tree_23 = a_in[23]^b_in[23];
endmodule // adder_tree_23
module adder_tree_24(
	input  [24:0] a_in,
	input  [24:0] b_in,
	input   n38_tree_30,
	input   n39_tree_30,
	input   n114_tree_28,
	output  sum
);
// adder_forest tree_24
	wire n97_tree_24, n103_tree_24;
    assign n97_tree_24 = (n114_tree_28&n39_tree_30)|n38_tree_30;
    assign sum = n97_tree_24^n103_tree_24;
    assign n103_tree_24 = a_in[24]^b_in[24];
endmodule // adder_tree_24
module adder_tree_25(
	input  [25:0] a_in,
	input  [25:0] b_in,
	input   n33_tree_32,
	input   n32_tree_32,
	input   n38_tree_30,
	input   n39_tree_30,
	input   n114_tree_28,
	output  sum
);
// adder_forest tree_25
	wire n3_tree_25, n100_tree_25, n101_tree_25, n107_tree_25;
    assign n100_tree_25 = n33_tree_32&n39_tree_30;
    assign n3_tree_25 = (n38_tree_30&n33_tree_32)|n32_tree_32;
    assign n101_tree_25 = (n114_tree_28&n100_tree_25)|n3_tree_25;
    assign sum = n101_tree_25^n107_tree_25;
    assign n107_tree_25 = a_in[25]^b_in[25];
endmodule // adder_tree_25
module adder_tree_26(
	input  [26:0] a_in,
	input  [26:0] b_in,
	input   n26_tree_32,
	input   n27_tree_32,
	input   n38_tree_30,
	input   n39_tree_30,
	input   n114_tree_28,
	output  sum
);
// adder_forest tree_26
	wire n6_tree_26, n7_tree_26, n105_tree_26, n111_tree_26;
    assign n7_tree_26 = n27_tree_32&n39_tree_30;
    assign n6_tree_26 = (n38_tree_30&n27_tree_32)|n26_tree_32;
    assign n105_tree_26 = (n114_tree_28&n7_tree_26)|n6_tree_26;
    assign sum = n105_tree_26^n111_tree_26;
    assign n111_tree_26 = a_in[26]^b_in[26];
endmodule // adder_tree_26
module adder_tree_27(
	input  [27:0] a_in,
	input  [27:0] b_in,
	input   n25_tree_32,
	input   n24_tree_32,
	input   n26_tree_32,
	input   n27_tree_32,
	input   n38_tree_30,
	input   n39_tree_30,
	input   n114_tree_28,
	output  sum
);
// adder_forest tree_27
	wire n3_tree_27, n10_tree_27, n11_tree_27, n108_tree_27, n109_tree_27, n115_tree_27;
    assign n108_tree_27 = n25_tree_32&n27_tree_32;
    assign n3_tree_27 = (n26_tree_32&n25_tree_32)|n24_tree_32;
    assign n11_tree_27 = n108_tree_27&n39_tree_30;
    assign n10_tree_27 = (n38_tree_30&n108_tree_27)|n3_tree_27;
    assign n109_tree_27 = (n114_tree_28&n11_tree_27)|n10_tree_27;
    assign sum = n109_tree_27^n115_tree_27;
    assign n115_tree_27 = a_in[27]^b_in[27];
endmodule // adder_tree_27
module adder_tree_28(
	input  [28:0] a_in,
	input  [28:0] b_in,
	input   n18_tree_31,
	input   n19_tree_31,
	input   n38_tree_30,
	input   n39_tree_30,
	input   n70_tree_30,
	input   n71_tree_30,
	input   n119_tree_29,
	output  sum,
	output  n114_tree_28
);
// adder_forest tree_28
	wire n14_tree_28, n15_tree_28, n113_tree_28, n119_tree_28;
    assign n15_tree_28 = n19_tree_31&n39_tree_30;
    assign n14_tree_28 = (n38_tree_30&n19_tree_31)|n18_tree_31;
    assign n113_tree_28 = (n114_tree_28&n15_tree_28)|n14_tree_28;
    assign n114_tree_28 = (n119_tree_29&n71_tree_30)|n70_tree_30;
    assign sum = n113_tree_28^n119_tree_28;
    assign n119_tree_28 = a_in[28]^b_in[28];
endmodule // adder_tree_28
module adder_tree_29(
	input  [29:0] a_in,
	input  [29:0] b_in,
	input   n17_tree_32,
	input   n16_tree_32,
	input   n18_tree_31,
	input   n19_tree_31,
	input   n38_tree_30,
	input   n39_tree_30,
	input   n70_tree_30,
	input   n71_tree_30,
	input   n98_tree_31,
	input   n99_tree_31,
	input   n124_tree_30,
	output  sum,
	output  n119_tree_29
);
// adder_forest tree_29
	wire n3_tree_29, n18_tree_29, n19_tree_29, n116_tree_29, n117_tree_29, n118_tree_29, n123_tree_29;
    assign n116_tree_29 = n17_tree_32&n19_tree_31;
    assign n3_tree_29 = (n18_tree_31&n17_tree_32)|n16_tree_32;
    assign n19_tree_29 = n116_tree_29&n39_tree_30;
    assign n18_tree_29 = (n38_tree_30&n116_tree_29)|n3_tree_29;
    assign n117_tree_29 = (n118_tree_29&n19_tree_29)|n18_tree_29;
    assign n118_tree_29 = (n119_tree_29&n71_tree_30)|n70_tree_30;
    assign n119_tree_29 = (n124_tree_30&n99_tree_31)|n98_tree_31;
    assign sum = n117_tree_29^n123_tree_29;
    assign n123_tree_29 = a_in[29]^b_in[29];
endmodule // adder_tree_29
module adder_tree_30(
	input  [30:0] a_in,
	input  [30:0] b_in,
	input   n10_tree_32,
	input   n11_tree_32,
	input   n18_tree_31,
	input   n19_tree_31,
	input   n34_tree_31,
	input   n35_tree_31,
	input   n50_tree_31,
	input   n51_tree_31,
	input   n66_tree_31,
	input   n67_tree_31,
	input   n82_tree_31,
	input   n83_tree_31,
	input   n98_tree_31,
	input   n99_tree_31,
	input   n114_tree_32,
	input   n115_tree_32,
	input   n129_tree_31,
	output  sum,
	output  n38_tree_30,
	output  n39_tree_30,
	output  n70_tree_30,
	output  n71_tree_30,
	output  n124_tree_30
);
// adder_forest tree_30
	wire n6_tree_30, n7_tree_30, n22_tree_30, n23_tree_30, n121_tree_30, n122_tree_30, n123_tree_30, n127_tree_30;
    assign n7_tree_30 = n11_tree_32&n19_tree_31;
    assign n6_tree_30 = (n18_tree_31&n11_tree_32)|n10_tree_32;
    assign n23_tree_30 = n7_tree_30&n39_tree_30;
    assign n22_tree_30 = (n38_tree_30&n7_tree_30)|n6_tree_30;
    assign n39_tree_30 = n35_tree_31&n51_tree_31;
    assign n38_tree_30 = (n50_tree_31&n35_tree_31)|n34_tree_31;
    assign n71_tree_30 = n67_tree_31&n83_tree_31;
    assign n70_tree_30 = (n82_tree_31&n67_tree_31)|n66_tree_31;
    assign n121_tree_30 = (n122_tree_30&n23_tree_30)|n22_tree_30;
    assign n122_tree_30 = (n123_tree_30&n71_tree_30)|n70_tree_30;
    assign n123_tree_30 = (n124_tree_30&n99_tree_31)|n98_tree_31;
    assign n124_tree_30 = (n129_tree_31&n115_tree_32)|n114_tree_32;
    assign sum = n121_tree_30^n127_tree_30;
    assign n127_tree_30 = a_in[30]^b_in[30];
endmodule // adder_tree_30
module adder_tree_31(
	input  [31:0] a_in,
	input  [31:0] b_in,
	input   n125_tree_32,
	input   n124_tree_32,
	input   n9_tree_32,
	input   n8_tree_32,
	input   n10_tree_32,
	input   n11_tree_32,
	input   n18_tree_32,
	input   n19_tree_32,
	input   n26_tree_32,
	input   n27_tree_32,
	input   n34_tree_32,
	input   n35_tree_32,
	input   n42_tree_32,
	input   n43_tree_32,
	input   n50_tree_32,
	input   n51_tree_32,
	input   n58_tree_32,
	input   n59_tree_32,
	input   n66_tree_32,
	input   n67_tree_32,
	input   n74_tree_32,
	input   n75_tree_32,
	input   n82_tree_32,
	input   n83_tree_32,
	input   n90_tree_32,
	input   n91_tree_32,
	input   n98_tree_32,
	input   n99_tree_32,
	input   n106_tree_32,
	input   n107_tree_32,
	input   n114_tree_32,
	input   n115_tree_32,
	input   n134_tree_32,
	output  sum,
	output  n18_tree_31,
	output  n19_tree_31,
	output  n34_tree_31,
	output  n35_tree_31,
	output  n50_tree_31,
	output  n51_tree_31,
	output  n66_tree_31,
	output  n67_tree_31,
	output  n82_tree_31,
	output  n83_tree_31,
	output  n98_tree_31,
	output  n99_tree_31,
	output  n129_tree_31
);
// adder_forest tree_31
	wire n3_tree_31, n10_tree_31, n11_tree_31, n26_tree_31, n27_tree_31, n42_tree_31, n43_tree_31, n74_tree_31, n75_tree_31, n124_tree_31, n125_tree_31, n126_tree_31, n127_tree_31, n128_tree_31, n131_tree_31;
    assign n124_tree_31 = n9_tree_32&n11_tree_32;
    assign n3_tree_31 = (n10_tree_32&n9_tree_32)|n8_tree_32;
    assign n11_tree_31 = n124_tree_31&n19_tree_31;
    assign n10_tree_31 = (n18_tree_31&n124_tree_31)|n3_tree_31;
    assign n19_tree_31 = n19_tree_32&n27_tree_32;
    assign n18_tree_31 = (n26_tree_32&n19_tree_32)|n18_tree_32;
    assign n27_tree_31 = n11_tree_31&n43_tree_31;
    assign n26_tree_31 = (n42_tree_31&n11_tree_31)|n10_tree_31;
    assign n35_tree_31 = n35_tree_32&n43_tree_32;
    assign n34_tree_31 = (n42_tree_32&n35_tree_32)|n34_tree_32;
    assign n43_tree_31 = n35_tree_31&n51_tree_31;
    assign n42_tree_31 = (n50_tree_31&n35_tree_31)|n34_tree_31;
    assign n51_tree_31 = n51_tree_32&n59_tree_32;
    assign n50_tree_31 = (n58_tree_32&n51_tree_32)|n50_tree_32;
    assign n67_tree_31 = n67_tree_32&n75_tree_32;
    assign n66_tree_31 = (n74_tree_32&n67_tree_32)|n66_tree_32;
    assign n75_tree_31 = n67_tree_31&n83_tree_31;
    assign n74_tree_31 = (n82_tree_31&n67_tree_31)|n66_tree_31;
    assign n83_tree_31 = n83_tree_32&n91_tree_32;
    assign n82_tree_31 = (n90_tree_32&n83_tree_32)|n82_tree_32;
    assign n99_tree_31 = n99_tree_32&n107_tree_32;
    assign n98_tree_31 = (n106_tree_32&n99_tree_32)|n98_tree_32;
    assign n125_tree_31 = (n126_tree_31&n27_tree_31)|n26_tree_31;
    assign n126_tree_31 = (n127_tree_31&n75_tree_31)|n74_tree_31;
    assign n127_tree_31 = (n128_tree_31&n99_tree_31)|n98_tree_31;
    assign n128_tree_31 = (n129_tree_31&n115_tree_32)|n114_tree_32;
    assign n129_tree_31 = (n134_tree_32&n125_tree_32)|n124_tree_32;
    assign sum = n125_tree_31^n131_tree_31;
    assign n131_tree_31 = a_in[31]^b_in[31];
endmodule // adder_tree_31
module adder_tree_32(
	input  [32:0] a_in,
	input  [32:0] b_in,
	output  sum,
	output  n125_tree_32,
	output  n124_tree_32,
	output  n121_tree_32,
	output  n120_tree_32,
	output  n117_tree_32,
	output  n116_tree_32,
	output  n113_tree_32,
	output  n112_tree_32,
	output  n109_tree_32,
	output  n108_tree_32,
	output  n105_tree_32,
	output  n104_tree_32,
	output  n101_tree_32,
	output  n100_tree_32,
	output  n97_tree_32,
	output  n96_tree_32,
	output  n93_tree_32,
	output  n92_tree_32,
	output  n89_tree_32,
	output  n88_tree_32,
	output  n85_tree_32,
	output  n84_tree_32,
	output  n81_tree_32,
	output  n80_tree_32,
	output  n77_tree_32,
	output  n76_tree_32,
	output  n73_tree_32,
	output  n72_tree_32,
	output  n69_tree_32,
	output  n68_tree_32,
	output  n65_tree_32,
	output  n64_tree_32,
	output  n61_tree_32,
	output  n60_tree_32,
	output  n57_tree_32,
	output  n56_tree_32,
	output  n53_tree_32,
	output  n52_tree_32,
	output  n49_tree_32,
	output  n48_tree_32,
	output  n45_tree_32,
	output  n44_tree_32,
	output  n41_tree_32,
	output  n40_tree_32,
	output  n37_tree_32,
	output  n36_tree_32,
	output  n33_tree_32,
	output  n32_tree_32,
	output  n29_tree_32,
	output  n28_tree_32,
	output  n25_tree_32,
	output  n24_tree_32,
	output  n21_tree_32,
	output  n20_tree_32,
	output  n17_tree_32,
	output  n16_tree_32,
	output  n13_tree_32,
	output  n12_tree_32,
	output  n9_tree_32,
	output  n8_tree_32,
	output  n10_tree_32,
	output  n11_tree_32,
	output  n18_tree_32,
	output  n19_tree_32,
	output  n26_tree_32,
	output  n27_tree_32,
	output  n34_tree_32,
	output  n35_tree_32,
	output  n42_tree_32,
	output  n43_tree_32,
	output  n50_tree_32,
	output  n51_tree_32,
	output  n58_tree_32,
	output  n59_tree_32,
	output  n66_tree_32,
	output  n67_tree_32,
	output  n74_tree_32,
	output  n75_tree_32,
	output  n82_tree_32,
	output  n83_tree_32,
	output  n90_tree_32,
	output  n91_tree_32,
	output  n98_tree_32,
	output  n99_tree_32,
	output  n106_tree_32,
	output  n107_tree_32,
	output  n114_tree_32,
	output  n115_tree_32,
	output  n134_tree_32
);
// adder_forest tree_32
	wire n3_tree_32, n4_tree_32, n5_tree_32, n6_tree_32, n7_tree_32, n14_tree_32, n15_tree_32, n22_tree_32, n23_tree_32, n30_tree_32, n31_tree_32, n38_tree_32, n39_tree_32, n46_tree_32, n47_tree_32, n54_tree_32, n55_tree_32, n70_tree_32, n71_tree_32, n78_tree_32, n79_tree_32, n86_tree_32, n87_tree_32, n102_tree_32, n103_tree_32, n128_tree_32, n129_tree_32, n130_tree_32, n131_tree_32, n132_tree_32, n133_tree_32, n135_tree_32;
    assign n125_tree_32 = a_in[1]^b_in[1];
    assign n124_tree_32 = a_in[1]&b_in[1];
    assign n121_tree_32 = a_in[2]^b_in[2];
    assign n120_tree_32 = a_in[2]&b_in[2];
    assign n117_tree_32 = a_in[3]^b_in[3];
    assign n116_tree_32 = a_in[3]&b_in[3];
    assign n113_tree_32 = a_in[4]^b_in[4];
    assign n112_tree_32 = a_in[4]&b_in[4];
    assign n109_tree_32 = a_in[5]^b_in[5];
    assign n108_tree_32 = a_in[5]&b_in[5];
    assign n105_tree_32 = a_in[6]^b_in[6];
    assign n104_tree_32 = a_in[6]&b_in[6];
    assign n101_tree_32 = a_in[7]^b_in[7];
    assign n100_tree_32 = a_in[7]&b_in[7];
    assign n97_tree_32 = a_in[8]^b_in[8];
    assign n96_tree_32 = a_in[8]&b_in[8];
    assign n93_tree_32 = a_in[9]^b_in[9];
    assign n92_tree_32 = a_in[9]&b_in[9];
    assign n89_tree_32 = a_in[10]^b_in[10];
    assign n88_tree_32 = a_in[10]&b_in[10];
    assign n85_tree_32 = a_in[11]^b_in[11];
    assign n84_tree_32 = a_in[11]&b_in[11];
    assign n81_tree_32 = a_in[12]^b_in[12];
    assign n80_tree_32 = a_in[12]&b_in[12];
    assign n77_tree_32 = a_in[13]^b_in[13];
    assign n76_tree_32 = a_in[13]&b_in[13];
    assign n73_tree_32 = a_in[14]^b_in[14];
    assign n72_tree_32 = a_in[14]&b_in[14];
    assign n69_tree_32 = a_in[15]^b_in[15];
    assign n68_tree_32 = a_in[15]&b_in[15];
    assign n65_tree_32 = a_in[16]^b_in[16];
    assign n64_tree_32 = a_in[16]&b_in[16];
    assign n61_tree_32 = a_in[17]^b_in[17];
    assign n60_tree_32 = a_in[17]&b_in[17];
    assign n57_tree_32 = a_in[18]^b_in[18];
    assign n56_tree_32 = a_in[18]&b_in[18];
    assign n53_tree_32 = a_in[19]^b_in[19];
    assign n52_tree_32 = a_in[19]&b_in[19];
    assign n49_tree_32 = a_in[20]^b_in[20];
    assign n48_tree_32 = a_in[20]&b_in[20];
    assign n45_tree_32 = a_in[21]^b_in[21];
    assign n44_tree_32 = a_in[21]&b_in[21];
    assign n41_tree_32 = a_in[22]^b_in[22];
    assign n40_tree_32 = a_in[22]&b_in[22];
    assign n37_tree_32 = a_in[23]^b_in[23];
    assign n36_tree_32 = a_in[23]&b_in[23];
    assign n33_tree_32 = a_in[24]^b_in[24];
    assign n32_tree_32 = a_in[24]&b_in[24];
    assign n29_tree_32 = a_in[25]^b_in[25];
    assign n28_tree_32 = a_in[25]&b_in[25];
    assign n25_tree_32 = a_in[26]^b_in[26];
    assign n24_tree_32 = a_in[26]&b_in[26];
    assign n21_tree_32 = a_in[27]^b_in[27];
    assign n20_tree_32 = a_in[27]&b_in[27];
    assign n17_tree_32 = a_in[28]^b_in[28];
    assign n16_tree_32 = a_in[28]&b_in[28];
    assign n13_tree_32 = a_in[29]^b_in[29];
    assign n12_tree_32 = a_in[29]&b_in[29];
    assign n9_tree_32 = a_in[30]^b_in[30];
    assign n8_tree_32 = a_in[30]&b_in[30];
    assign n5_tree_32 = a_in[31]^b_in[31];
    assign n4_tree_32 = a_in[31]&b_in[31];
    assign n128_tree_32 = n5_tree_32&n9_tree_32;
    assign n3_tree_32 = (n8_tree_32&n5_tree_32)|n4_tree_32;
    assign n7_tree_32 = n128_tree_32&n11_tree_32;
    assign n6_tree_32 = (n10_tree_32&n128_tree_32)|n3_tree_32;
    assign n11_tree_32 = n13_tree_32&n17_tree_32;
    assign n10_tree_32 = (n16_tree_32&n13_tree_32)|n12_tree_32;
    assign n15_tree_32 = n7_tree_32&n23_tree_32;
    assign n14_tree_32 = (n22_tree_32&n7_tree_32)|n6_tree_32;
    assign n19_tree_32 = n21_tree_32&n25_tree_32;
    assign n18_tree_32 = (n24_tree_32&n21_tree_32)|n20_tree_32;
    assign n23_tree_32 = n19_tree_32&n27_tree_32;
    assign n22_tree_32 = (n26_tree_32&n19_tree_32)|n18_tree_32;
    assign n27_tree_32 = n29_tree_32&n33_tree_32;
    assign n26_tree_32 = (n32_tree_32&n29_tree_32)|n28_tree_32;
    assign n31_tree_32 = n15_tree_32&n47_tree_32;
    assign n30_tree_32 = (n46_tree_32&n15_tree_32)|n14_tree_32;
    assign n35_tree_32 = n37_tree_32&n41_tree_32;
    assign n34_tree_32 = (n40_tree_32&n37_tree_32)|n36_tree_32;
    assign n39_tree_32 = n35_tree_32&n43_tree_32;
    assign n38_tree_32 = (n42_tree_32&n35_tree_32)|n34_tree_32;
    assign n43_tree_32 = n45_tree_32&n49_tree_32;
    assign n42_tree_32 = (n48_tree_32&n45_tree_32)|n44_tree_32;
    assign n47_tree_32 = n39_tree_32&n55_tree_32;
    assign n46_tree_32 = (n54_tree_32&n39_tree_32)|n38_tree_32;
    assign n51_tree_32 = n53_tree_32&n57_tree_32;
    assign n50_tree_32 = (n56_tree_32&n53_tree_32)|n52_tree_32;
    assign n55_tree_32 = n51_tree_32&n59_tree_32;
    assign n54_tree_32 = (n58_tree_32&n51_tree_32)|n50_tree_32;
    assign n59_tree_32 = n61_tree_32&n65_tree_32;
    assign n58_tree_32 = (n64_tree_32&n61_tree_32)|n60_tree_32;
    assign n67_tree_32 = n69_tree_32&n73_tree_32;
    assign n66_tree_32 = (n72_tree_32&n69_tree_32)|n68_tree_32;
    assign n71_tree_32 = n67_tree_32&n75_tree_32;
    assign n70_tree_32 = (n74_tree_32&n67_tree_32)|n66_tree_32;
    assign n75_tree_32 = n77_tree_32&n81_tree_32;
    assign n74_tree_32 = (n80_tree_32&n77_tree_32)|n76_tree_32;
    assign n79_tree_32 = n71_tree_32&n87_tree_32;
    assign n78_tree_32 = (n86_tree_32&n71_tree_32)|n70_tree_32;
    assign n83_tree_32 = n85_tree_32&n89_tree_32;
    assign n82_tree_32 = (n88_tree_32&n85_tree_32)|n84_tree_32;
    assign n87_tree_32 = n83_tree_32&n91_tree_32;
    assign n86_tree_32 = (n90_tree_32&n83_tree_32)|n82_tree_32;
    assign n91_tree_32 = n93_tree_32&n97_tree_32;
    assign n90_tree_32 = (n96_tree_32&n93_tree_32)|n92_tree_32;
    assign n99_tree_32 = n101_tree_32&n105_tree_32;
    assign n98_tree_32 = (n104_tree_32&n101_tree_32)|n100_tree_32;
    assign n103_tree_32 = n99_tree_32&n107_tree_32;
    assign n102_tree_32 = (n106_tree_32&n99_tree_32)|n98_tree_32;
    assign n107_tree_32 = n109_tree_32&n113_tree_32;
    assign n106_tree_32 = (n112_tree_32&n109_tree_32)|n108_tree_32;
    assign n115_tree_32 = n117_tree_32&n121_tree_32;
    assign n114_tree_32 = (n120_tree_32&n117_tree_32)|n116_tree_32;
    assign n129_tree_32 = (n130_tree_32&n31_tree_32)|n30_tree_32;
    assign n130_tree_32 = (n131_tree_32&n79_tree_32)|n78_tree_32;
    assign n131_tree_32 = (n132_tree_32&n103_tree_32)|n102_tree_32;
    assign n132_tree_32 = (n133_tree_32&n115_tree_32)|n114_tree_32;
    assign n133_tree_32 = (n134_tree_32&n125_tree_32)|n124_tree_32;
    assign n134_tree_32 = a_in[0]&b_in[0];
    assign sum = n129_tree_32^n135_tree_32;
    assign n135_tree_32 = a_in[32]^b_in[32];
endmodule // adder_tree_32
`endif