// wishbone.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module wishbone#(
    parameter SLAVE_SAYISI = 1
)(
);

endmodule