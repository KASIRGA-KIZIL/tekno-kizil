@40000000
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00
@40000048
93 00 00 00 93 01 00 00 13 02 00 00 93 02 00 00
13 03 00 00 93 03 00 00 13 04 00 00 93 04 00 00
13 05 00 00 93 05 00 00 13 06 00 00 93 06 00 00
13 07 00 00 93 07 00 00 13 08 00 00 93 08 00 00
13 09 00 00 93 09 00 00 13 0A 00 00 93 0A 00 00
13 0B 00 00 93 0B 00 00 13 0C 00 00 93 0C 00 00
13 0D 00 00 93 0D 00 00 13 0E 00 00 93 0E 00 00
13 0F 00 00 93 0F 00 00 97 41 00 00 93 81 01 03
17 72 00 00 13 02 F2 E2 13 72 02 FC 13 05 00 00
93 05 10 00 63 70 B5 00 13 01 15 00 13 11 E1 00
33 01 41 00 13 16 E5 00 33 02 C2 00 EF 20 10 64
6F 00 00 00 33 67 B5 00 93 03 F0 FF 13 77 37 00
63 10 07 10 B7 87 7F 7F 93 87 F7 F7 03 26 05 00
83 A6 05 00 B3 72 F6 00 33 63 F6 00 B3 82 F2 00
B3 E2 62 00 63 92 72 10 63 16 D6 08 03 26 45 00
83 A6 45 00 B3 72 F6 00 33 63 F6 00 B3 82 F2 00
B3 E2 62 00 63 9E 72 0C 63 16 D6 06 03 26 85 00
83 A6 85 00 B3 72 F6 00 33 63 F6 00 B3 82 F2 00
B3 E2 62 00 63 98 72 0C 63 16 D6 04 03 26 C5 00
83 A6 C5 00 B3 72 F6 00 33 63 F6 00 B3 82 F2 00
B3 E2 62 00 63 92 72 0C 63 16 D6 02 03 26 05 01
83 A6 05 01 B3 72 F6 00 33 63 F6 00 B3 82 F2 00
B3 E2 62 00 63 9C 72 0A 13 05 45 01 93 85 45 01
E3 0E D6 F4 13 17 06 01 93 97 06 01 63 1E F7 00
13 57 06 01 93 D7 06 01 33 05 F7 40 93 75 F5 0F
63 90 05 02 67 80 00 00 13 57 07 01 93 D7 07 01
33 05 F7 40 93 75 F5 0F 63 94 05 00 67 80 00 00
13 77 F7 0F 93 F7 F7 0F 33 05 F7 40 67 80 00 00
03 46 05 00 83 C6 05 00 13 05 15 00 93 85 15 00
63 14 D6 00 E3 16 06 FE 33 05 D6 40 67 80 00 00
13 05 45 00 93 85 45 00 E3 1C D6 FC 13 05 00 00
67 80 00 00 13 05 85 00 93 85 85 00 E3 12 D6 FC
13 05 00 00 67 80 00 00 13 05 C5 00 93 85 C5 00
E3 18 D6 FA 13 05 00 00 67 80 00 00 13 05 05 01
93 85 05 01 E3 1E D6 F8 13 05 00 00 67 80 00 00
13 01 01 FD 23 26 71 01 93 0B 06 00 13 D6 45 01
23 24 81 02 23 20 21 03 23 2E 31 01 23 28 61 01
13 94 C5 00 23 26 11 02 23 22 91 02 23 2C 41 01
23 2A 51 01 13 76 F6 7F 13 0B 05 00 13 89 06 00
13 54 C4 00 93 D9 F5 01 63 0E 06 08 93 07 F0 7F
63 0E F6 0E 93 56 D5 01 13 14 34 00 B3 E6 86 00
B7 07 80 00 33 EA F6 00 93 14 35 00 93 0A 16 C0
13 0B 00 00 93 57 49 01 13 14 C9 00 93 F7 F7 7F
13 54 C4 00 13 59 F9 01 63 80 07 10 13 07 F0 7F
63 84 E7 16 13 14 34 00 13 D7 DB 01 33 67 87 00
37 04 80 00 33 64 87 00 13 9F 3B 00 93 86 17 C0
93 05 00 00 93 17 2B 00 B3 E7 B7 00 33 86 DA 40
93 87 F7 FF 93 06 E0 00 33 C7 29 01 63 EA F6 18
93 97 27 00 93 86 01 04 B3 87 D7 00 83 A7 07 00
67 80 07 00 33 6A A4 00 63 00 0A 08 63 0E 04 02
13 05 04 00 EF 00 50 63 93 07 55 FF 93 06 D0 01
13 07 85 FF B3 86 F6 40 33 14 E4 00 B3 56 DB 00
33 EA 86 00 33 14 EB 00 13 06 D0 C0 B3 0A A6 40
93 04 04 00 6F F0 DF F4 EF 00 10 60 13 0A 05 00
93 07 5A 01 13 07 C0 01 13 05 05 02 E3 50 F7 FC
13 0A 8A FF 33 1A 4B 01 6F F0 1F FD 33 6A A4 00
63 04 0A 02 93 04 05 00 13 0A 04 00 93 0A F0 7F
13 0B 30 00 6F F0 1F F1 93 04 00 00 93 0A 00 00
13 0B 10 00 6F F0 1F F0 93 04 00 00 93 0A F0 7F
13 0B 20 00 6F F0 1F EF 33 6F 74 01 63 02 0F 08
63 00 04 04 13 05 04 00 EF 00 10 59 13 07 55 FF
93 07 D0 01 93 06 85 FF B3 87 E7 40 33 14 D4 00
B3 D7 FB 00 B3 E7 87 00 33 94 DB 00 93 06 D0 C0
13 0F 04 00 B3 86 A6 40 13 84 07 00 6F F0 5F EE
13 85 0B 00 EF 00 50 55 93 07 05 00 13 87 57 01
93 06 C0 01 13 05 05 02 E3 DC E6 FA 93 87 87 FF
B3 97 FB 00 6F F0 9F FC 33 6F 74 01 63 02 0F 02
13 8F 0B 00 93 06 F0 7F 93 05 30 00 6F F0 9F EA
13 04 00 00 93 06 00 00 93 05 10 00 6F F0 9F E9
13 04 00 00 93 06 F0 7F 93 05 20 00 6F F0 9F E8
13 87 09 00 13 04 0A 00 13 8F 04 00 93 07 20 00
63 02 FB 46 93 07 30 00 63 04 FB 44 93 07 10 00
63 12 FB 2C 13 04 00 00 93 06 00 00 6F 00 80 3F
63 66 44 01 63 1E 8A 34 63 EC E4 35 93 16 FA 01
93 D7 14 00 13 93 F4 01 13 5A 1A 00 B3 E4 F6 00
13 14 84 00 93 58 04 01 B3 5E 1A 03 93 55 8F 01
B3 E5 85 00 13 98 05 01 13 58 08 01 93 D7 04 01
13 15 8F 00 B3 76 1A 03 33 0E D8 03 93 96 06 01
B3 E7 D7 00 93 86 0E 00 63 FE C7 01 B3 87 F5 00
93 86 FE FF 63 E8 B7 00 63 F6 C7 01 93 86 EE FF
B3 87 B7 00 B3 87 C7 41 B3 DE 17 03 93 94 04 01
93 D4 04 01 B3 F7 17 03 33 0E D8 03 93 97 07 01
B3 E4 F4 00 93 87 0E 00 63 FE C4 01 B3 84 95 00
93 87 FE FF 63 E8 B4 00 63 F6 C4 01 93 87 EE FF
B3 84 B4 00 93 96 06 01 B7 03 01 00 B3 EF F6 00
B3 84 C4 41 13 8E F3 FF B3 F7 CF 01 13 DF 0F 01
93 5E 05 01 33 7E C5 01 B3 02 FE 02 33 04 CF 03
93 D6 02 01 B3 87 FE 02 B3 87 87 00 B3 86 F6 00
33 0F DF 03 63 F4 86 00 33 0F 7F 00 93 D7 06 01
B3 87 E7 01 37 0F 01 00 13 0F FF FF B3 F6 E6 01
93 96 06 01 B3 F2 E2 01 B3 86 56 00 63 E8 F4 00
13 84 0F 00 63 98 F4 04 63 76 D3 04 33 0F A3 00
B3 32 6F 00 B3 83 B2 00 B3 84 74 00 13 84 FF FF
13 03 0F 00 63 E6 95 00 63 96 95 02 63 94 02 02
63 E6 F4 00 63 90 97 02 63 7E DF 00 33 0F E5 01
13 03 0F 00 33 3F AF 00 33 0F BF 00 13 84 EF FF
B3 84 E4 01 B3 06 D3 40 B3 84 F4 40 33 33 D3 00
B3 84 64 40 13 0F F0 FF 63 86 95 12 B3 DF 14 03
93 D7 06 01 B3 F4 14 03 13 83 0F 00 33 0F F8 03
93 94 04 01 B3 E7 97 00 63 FE E7 01 B3 87 F5 00
13 83 FF FF 63 E8 B7 00 63 F6 E7 01 13 83 EF FF
B3 87 B7 00 B3 87 E7 41 33 DF 17 03 93 96 06 01
93 D6 06 01 B3 F7 17 03 33 08 E8 03 93 97 07 01
B3 E7 F6 00 93 06 0F 00 63 FE 07 01 B3 87 F5 00
93 06 FF FF 63 E8 B7 00 63 F6 07 01 93 06 EF FF
B3 87 B7 00 13 13 03 01 33 63 D3 00 93 16 03 01
93 D6 06 01 93 58 03 01 33 8F C6 03 B3 87 07 41
33 8E C8 03 B3 88 1E 03 B3 8E DE 02 93 56 0F 01
B3 8E CE 01 B3 86 D6 01 63 F6 C6 01 37 08 01 00
B3 88 08 01 13 D8 06 01 33 08 18 01 B7 08 01 00
93 88 F8 FF B3 F6 16 01 93 96 06 01 33 7F 1F 01
B3 86 E6 01 63 E8 07 01 13 0F 03 00 63 92 07 05
63 82 06 04 B3 87 F5 00 13 0F F3 FF 93 88 07 00
63 E4 B7 02 63 E6 07 01 63 94 07 03 63 70 D5 02
13 0F E3 FF 13 13 15 00 B3 38 A3 00 B3 88 B8 00
B3 88 17 01 13 05 03 00 63 94 08 01 63 84 A6 00
13 6F 1F 00 93 07 F6 3F 63 50 F0 0C 93 76 7F 00
63 80 06 02 93 76 FF 00 93 05 40 00 63 8A B6 00
93 06 4F 00 B3 B5 E6 01 33 04 B4 00 13 8F 06 00
B7 06 00 01 B3 76 D4 00 63 8A 06 00 B7 07 00 FF
93 87 F7 FF 33 74 F4 00 93 07 06 40 93 06 E0 7F
63 C2 F6 14 93 16 D4 01 13 5F 3F 00 B3 E6 E6 01
13 54 34 00 13 14 C4 00 13 54 C4 00 93 97 47 01
83 20 C1 02 B3 E7 87 00 03 24 81 02 13 17 F7 01
33 E6 E7 00 83 24 41 02 03 29 01 02 83 29 C1 01
03 2A 81 01 83 2A 41 01 03 2B 01 01 83 2B C1 00
13 85 06 00 93 05 06 00 13 01 01 03 67 80 00 00
13 06 F6 FF 13 03 00 00 6F F0 9F CB 13 07 09 00
13 8B 05 00 6F F0 9F C6 93 05 10 00 63 8C 07 00
B3 85 F5 40 93 06 80 03 E3 C6 B6 C6 93 06 F0 01
63 C6 B6 06 13 06 E6 41 B3 57 BF 00 33 1F CF 00
33 3F E0 01 33 16 C4 00 33 6F CF 00 B3 E7 E7 01
33 54 B4 00 93 F6 77 00 63 80 06 02 93 F6 F7 00
13 06 40 00 63 8A C6 00 93 86 47 00 33 B6 F6 00
33 04 C4 00 93 87 06 00 B7 06 80 00 B3 76 D4 00
63 9A 06 06 93 16 D4 01 93 D7 37 00 B3 E6 F6 00
13 54 34 00 93 07 00 00 6F F0 DF F1 93 06 10 FE
B3 87 F6 40 13 05 00 02 B3 57 F4 00 93 06 00 00
63 86 A5 00 13 06 E6 43 B3 16 C4 00 B3 E6 E6 01
B3 36 D0 00 B3 E7 D7 00 13 04 00 00 6F F0 9F F8
37 04 08 00 93 06 00 00 93 07 F0 7F 13 07 00 00
6F F0 5F ED 13 04 00 00 93 06 00 00 93 07 F0 7F
6F F0 5F EC 13 04 00 00 93 06 00 00 93 07 10 00
6F F0 5F EB 13 01 01 FF 23 24 81 00 23 26 11 00
13 04 05 00 63 02 05 06 EF 00 10 05 13 07 E0 41
93 07 A0 00 33 07 A7 40 63 C0 A7 04 93 07 B0 00
B3 87 A7 40 13 05 55 01 B3 57 F4 00 33 14 A4 00
83 20 C1 00 13 05 04 00 93 97 C7 00 03 24 81 00
13 17 47 01 93 D7 C7 00 B3 66 F7 00 93 85 06 00
13 01 01 01 67 80 00 00 13 05 55 FF B3 17 A4 00
13 04 00 00 6F F0 DF FC 93 07 00 00 13 07 00 00
6F F0 1F FC 13 01 01 FE 23 2A 91 00 93 54 75 01
23 28 21 01 23 26 31 01 23 24 41 01 13 17 95 00
23 2E 11 00 23 2C 81 00 23 22 51 01 93 F4 F4 0F
13 8A 05 00 93 59 97 00 13 59 F5 01 63 82 04 08
93 07 F0 0F 63 8E F4 08 13 97 39 00 B7 07 00 04
B3 69 F7 00 93 84 14 F8 93 0A 00 00 93 57 7A 01
13 14 9A 00 93 F7 F7 0F 13 54 94 00 13 5A FA 01
63 88 07 08 13 07 F0 0F 63 84 E7 0A 13 14 34 00
37 07 00 04 33 64 E4 00 93 87 17 F8 93 06 00 00
B3 84 F4 40 93 97 2A 00 B3 E7 D7 00 93 87 F7 FF
13 07 E0 00 33 46 49 01 63 64 F7 0C 93 97 27 00
13 87 C1 07 B3 87 E7 00 83 A7 07 00 67 80 07 00
63 8A 09 02 13 85 09 00 EF 00 00 72 93 07 B5 FF
93 04 A0 F8 B3 99 F9 00 B3 84 A4 40 6F F0 DF F7
93 04 F0 0F 93 0A 30 00 E3 9A 09 F6 93 0A 20 00
6F F0 DF F6 93 04 00 00 93 0A 10 00 6F F0 1F F6
63 0A 04 02 13 05 04 00 EF 00 00 6E 93 07 B5 FF
33 14 F4 00 93 07 A0 F8 B3 87 A7 40 6F F0 1F F7
93 07 F0 0F 93 06 30 00 E3 14 04 F6 93 06 20 00
6F F0 1F F6 93 07 00 00 93 06 10 00 6F F0 5F F5
13 06 09 00 13 84 09 00 93 86 0A 00 93 07 20 00
63 8A F6 1C 93 07 30 00 63 8E F6 1A 93 07 10 00
63 9C F6 0A 93 07 00 00 13 07 00 00 6F 00 40 0F
93 15 54 00 63 F4 89 12 93 84 F4 FF 93 07 00 00
13 D5 05 01 B3 D8 A9 02 B7 06 01 00 93 86 F6 FF
B3 F6 D5 00 93 D7 07 01 33 F7 A9 02 13 84 08 00
33 88 16 03 13 17 07 01 B3 E7 E7 00 63 FE 07 01
B3 87 F5 00 13 84 F8 FF 63 E8 B7 00 63 F6 07 01
13 84 E8 FF B3 87 B7 00 B3 87 07 41 33 D8 A7 02
B3 F7 A7 02 33 87 06 03 93 97 07 01 93 06 08 00
63 F2 E7 02 33 85 B7 00 B3 38 F5 00 93 06 F8 FF
93 07 05 00 63 98 08 00 63 76 E5 00 93 06 E8 FF
B3 07 B5 00 13 14 04 01 B3 87 E7 40 33 64 D4 00
B3 37 F0 00 33 64 F4 00 13 87 F4 07 63 5A E0 08
93 77 74 00 63 8A 07 00 93 77 F4 00 93 06 40 00
63 84 D7 00 13 04 44 00 B7 07 00 08 B3 77 F4 00
63 8A 07 00 B7 07 00 F8 93 87 F7 FF 33 74 F4 00
13 87 04 08 93 07 E0 0F 63 C6 E7 0C 93 57 34 00
83 20 C1 01 03 24 81 01 93 97 97 00 13 17 77 01
93 D7 97 00 33 67 F7 00 13 15 F6 01 83 24 41 01
03 29 01 01 83 29 C1 00 03 2A 81 00 83 2A 41 00
33 65 A7 00 13 01 01 02 67 80 00 00 93 97 F9 01
93 D9 19 00 6F F0 DF ED 13 06 0A 00 6F F0 1F EA
93 06 10 00 63 0C 07 00 B3 86 E6 40 93 05 B0 01
93 07 00 00 13 07 00 00 E3 CC D5 F8 93 84 E4 09
B3 56 D4 00 33 14 94 00 33 34 80 00 B3 E7 86 00
13 F7 77 00 63 0A 07 00 13 F7 F7 00 93 06 40 00
63 04 D7 00 93 87 47 00 37 07 00 04 33 F7 E7 00
93 D7 37 00 E3 0E 07 F4 93 07 00 00 13 07 10 00
6F F0 1F F5 B7 07 40 00 13 07 F0 0F 13 06 00 00
6F F0 1F F4 93 07 00 00 13 07 F0 0F 6F F0 5F F3
13 01 01 FE 23 28 21 01 13 59 75 01 23 2A 91 00
23 26 31 01 23 22 51 01 93 14 95 00 23 2E 11 00
23 2C 81 00 23 24 41 01 13 79 F9 0F 93 8A 05 00
93 D4 94 00 93 59 F5 01 63 06 09 18 93 07 F0 0F
63 02 F9 1A 93 94 34 00 B7 07 00 04 B3 E4 F4 00
13 09 19 F8 13 0A 00 00 93 D7 7A 01 13 94 9A 00
93 F7 F7 0F 13 54 94 00 93 DA FA 01 63 8C 07 18
13 07 F0 0F 63 88 E7 1A 13 14 34 00 37 07 00 04
33 64 E4 00 93 87 17 F8 13 07 00 00 33 09 F9 00
93 17 2A 00 B3 E7 E7 00 93 06 A0 00 33 C5 59 01
13 06 19 00 63 C4 F6 1E 93 06 20 00 63 CC F6 18
93 87 F7 FF 93 06 10 00 63 F8 F6 1A B7 08 01 00
13 88 F8 FF 13 D7 04 01 93 57 04 01 B3 76 04 01
B3 F4 04 01 B3 85 96 02 B3 06 D7 02 13 D4 05 01
33 07 F7 02 B3 87 97 02 B3 87 D7 00 33 04 F4 00
63 74 D4 00 33 07 17 01 B3 77 04 01 93 97 07 01
B3 F5 05 01 B3 87 B7 00 93 96 67 00 13 54 04 01
B3 36 D0 00 93 D7 A7 01 33 04 E4 00 B3 E7 F6 00
13 14 64 00 33 64 F4 00 B7 07 00 08 B3 77 F4 00
63 8E 07 16 93 57 14 00 13 74 14 00 33 E4 87 00
13 07 F6 07 63 58 E0 16 93 77 74 00 63 8A 07 00
93 77 F4 00 93 06 40 00 63 84 D7 00 13 04 44 00
B7 07 00 08 B3 77 F4 00 63 8A 07 00 B7 07 00 F8
93 87 F7 FF 33 74 F4 00 13 07 06 08 93 07 E0 0F
63 C4 E7 1A 93 57 34 00 83 20 C1 01 03 24 81 01
93 97 97 00 13 17 77 01 93 D7 97 00 33 67 F7 00
13 15 F5 01 83 24 41 01 03 29 01 01 83 29 C1 00
03 2A 81 00 83 2A 41 00 33 65 A7 00 13 01 01 02
67 80 00 00 63 8A 04 02 13 85 04 00 EF 00 C0 2E
93 07 B5 FF 13 09 A0 F8 B3 94 F4 00 33 09 A9 40
6F F0 5F E7 13 09 F0 0F 13 0A 30 00 E3 96 04 E6
13 0A 20 00 6F F0 5F E6 13 09 00 00 13 0A 10 00
6F F0 9F E5 63 0A 04 02 13 05 04 00 EF 00 C0 2A
93 07 B5 FF 33 14 F4 00 93 07 A0 F8 B3 87 A7 40
6F F0 9F E6 93 07 F0 0F 13 07 30 00 E3 10 04 E6
13 07 20 00 6F F0 9F E5 93 07 00 00 13 07 10 00
6F F0 DF E4 93 06 10 00 B3 97 F6 00 93 F6 07 53
63 98 06 04 93 F6 07 24 63 90 06 0C 93 F7 87 08
E3 8E 07 E4 13 85 0A 00 93 07 20 00 63 0E F7 0A
93 07 30 00 63 02 F7 0A 93 07 10 00 E3 12 F7 EC
93 07 00 00 13 07 00 00 6F F0 1F F0 93 06 F0 00
63 84 D7 08 93 06 B0 00 13 85 09 00 E3 84 D7 FC
13 84 04 00 13 07 0A 00 6F F0 1F FC 13 06 09 00
6F F0 1F E9 93 06 10 00 63 0C 07 00 B3 86 E6 40
93 05 B0 01 93 07 00 00 13 07 00 00 E3 CE D5 EA
13 06 E6 09 B3 56 D4 00 33 14 C4 00 33 34 80 00
B3 E7 86 00 13 F7 77 00 63 0A 07 00 13 F7 F7 00
93 06 40 00 63 04 D7 00 93 87 47 00 37 07 00 04
33 F7 E7 00 93 D7 37 00 E3 00 07 E8 93 07 00 00
13 07 10 00 6F F0 5F E7 B7 07 40 00 13 07 F0 0F
13 05 00 00 6F F0 5F E6 93 07 00 00 13 07 F0 0F
6F F0 9F E5 37 06 80 00 13 57 75 01 93 07 F6 FF
13 77 F7 0F 93 05 E0 07 B3 F7 A7 00 93 56 F5 01
63 D6 E5 04 93 05 D0 09 63 DA E5 00 37 05 00 80
13 45 F5 FF 33 85 A6 00 67 80 00 00 33 E5 C7 00
93 07 50 09 63 DC E7 00 13 07 A7 F6 33 15 E5 00
63 80 06 02 33 05 A0 40 67 80 00 00 93 07 60 09
B3 87 E7 40 33 55 F5 00 6F F0 9F FE 13 05 00 00
67 80 00 00 13 01 01 FF 23 26 11 00 23 24 81 00
23 22 91 00 93 07 05 00 63 06 05 0E 13 57 F5 41
33 44 A7 00 33 04 E4 40 93 54 F5 01 13 05 04 00
EF 00 80 0E 93 07 E0 09 B3 87 A7 40 13 07 60 09
63 40 F7 04 13 07 80 00 63 04 E5 0C 13 05 85 FF
33 14 A4 00 13 14 94 00 13 54 94 00 93 97 77 01
83 20 C1 00 B3 E7 87 00 03 24 81 00 13 95 F4 01
33 E5 A7 00 83 24 41 00 13 01 01 01 67 80 00 00
13 07 90 09 63 56 F7 06 13 07 50 00 33 07 A7 40
93 06 B5 01 33 57 E4 00 33 14 D4 00 33 34 80 00
33 64 87 00 37 07 00 FC 13 07 F7 FF 93 76 74 00
33 77 E4 00 63 8A 06 00 13 74 F4 00 93 06 40 00
63 04 D4 00 13 07 47 00 B7 06 00 04 B3 76 D7 00
63 8C 06 00 B7 07 00 FC 93 87 F7 FF 33 77 F7 00
93 07 F0 09 B3 87 A7 40 13 54 37 00 6F F0 9F F6
93 06 50 00 13 07 B5 FF E3 06 D5 FA 33 14 E4 00
6F F0 5F FA 93 04 00 00 13 04 00 00 6F F0 9F F4
93 07 60 09 6F F0 1F F4 B7 07 01 00 63 78 F5 02
93 37 05 10 93 C7 17 00 93 97 37 00 93 06 00 02
B3 86 F6 40 33 55 F5 00 93 87 81 0B B3 87 A7 00
03 C5 07 00 33 85 A6 40 67 80 00 00 37 07 00 01
93 07 00 01 E3 6C E5 FC 93 07 80 01 6F F0 1F FD
@400011E8
13 01 01 FA 23 2E 81 04 23 2C 91 04 93 F8 07 04
13 08 05 00 17 2F 00 00 13 0F CF 72 63 96 08 00
17 2F 00 00 13 0F 8F 6F 93 F2 07 01 63 98 02 44
13 F5 17 00 93 F4 17 01 93 0F 00 03 63 04 05 44
13 F5 27 00 93 F3 07 02 63 06 05 42 63 C6 05 44
13 F5 47 00 63 16 05 48 93 F7 87 00 13 04 00 00
63 86 07 00 93 86 F6 FF 13 04 00 02 63 8C 03 00
93 07 00 01 63 06 F6 4A 93 07 86 FF 93 B7 17 00
B3 86 F6 40 63 92 05 42 93 07 00 03 23 06 F1 00
13 05 10 00 13 03 C1 00 13 0E 05 00 63 54 E5 00
13 0E 07 00 B3 86 C6 41 63 90 04 0E 93 8E F6 FF
63 5A D0 48 33 07 00 41 93 08 50 00 93 77 37 00
63 FE D8 49 13 0F 08 00 63 80 07 04 93 08 00 02
23 00 18 01 13 77 27 00 13 0F 18 00 93 8E E6 FF
63 04 07 02 13 07 F8 FF A3 00 18 01 13 77 37 00
13 0F 28 00 93 8E D6 FF 63 18 07 00 13 0F 38 00
23 01 18 01 93 8E C6 FF B3 84 F6 40 93 F8 C4 FF
B3 07 F8 00 37 27 20 20 B3 88 F8 00 13 07 07 02
23 A0 E7 00 93 87 47 00 E3 9C F8 FE 13 F7 C4 FF
93 F4 34 00 B3 07 EF 00 B3 8E EE 40 63 82 04 04
13 07 00 02 23 80 E7 00 63 5C D0 03 A3 80 E7 00
93 08 10 00 63 86 1E 03 23 81 E7 00 93 08 20 00
63 80 1E 03 A3 81 E7 00 93 08 30 00 63 8A 1E 01
23 82 E7 00 93 08 40 00 63 84 1E 01 A3 82 E7 00
33 08 D8 00 93 06 F0 FF 63 06 04 00 23 00 88 00
13 08 18 00 63 8A 03 00 93 07 80 00 63 0A F6 36
93 07 00 01 63 04 F6 34 63 94 02 0E 93 88 F6 FF
63 5E D0 38 33 07 00 41 13 06 50 00 93 77 37 00
63 7A 16 39 93 0E 08 00 63 8E 07 02 23 00 F8 01
13 77 27 00 93 0E 18 00 93 88 E6 FF 63 04 07 02
13 07 F8 FF A3 00 F8 01 13 77 37 00 93 0E 28 00
93 88 D6 FF 63 18 07 00 93 0E 38 00 23 01 F8 01
93 88 C6 FF 13 97 8F 00 33 8F F6 40 13 96 0F 01
33 E7 EF 00 33 67 C7 00 93 92 8F 01 B3 07 F8 00
13 76 CF FF 33 67 57 00 33 06 F6 00 23 A0 E7 00
93 87 47 00 E3 9C C7 FE 13 77 CF FF 13 7F 3F 00
B3 87 EE 00 B3 88 E8 40 63 00 0F 04 23 80 F7 01
63 5C 10 03 A3 80 F7 01 13 07 10 00 63 86 E8 02
23 81 F7 01 13 07 20 00 63 80 E8 02 A3 81 F7 01
13 07 30 00 63 8A E8 00 23 82 F7 01 13 07 40 00
63 84 E8 00 A3 82 F7 01 33 08 D8 00 93 06 F0 FF
93 08 FE FF 63 5E C5 0D 33 0F AE 40 33 07 00 41
93 0E FF FF 13 06 50 00 93 77 37 00 63 78 D6 29
93 0E 08 00 63 80 07 04 13 06 00 03 23 00 C8 00
13 77 27 00 93 0E 18 00 93 08 EE FF 63 04 07 02
13 07 F8 FF A3 00 C8 00 13 77 37 00 93 0E 28 00
93 08 DE FF 63 18 07 00 93 0E 38 00 23 01 C8 00
93 08 CE FF 33 0E FF 40 13 76 CE FF B3 07 F8 00
37 37 30 30 33 06 F6 00 13 07 07 03 23 A0 E7 00
93 87 47 00 E3 1C F6 FE 93 77 3E 00 63 88 07 04
13 7E CE FF B3 87 CE 01 B3 88 C8 41 13 07 00 03
23 80 E7 00 13 86 F8 FF 63 5A 15 03 A3 80 E7 00
13 8E E8 FF 63 54 C5 02 23 81 E7 00 13 86 D8 FF
63 5E C5 01 A3 81 E7 00 93 88 C8 FF 63 58 C5 00
23 82 E7 00 63 54 15 01 A3 82 E7 00 33 08 E8 01
B3 07 B3 00 13 07 08 00 03 C5 07 00 13 86 07 00
13 07 17 00 A3 0F A7 FE 93 87 F7 FF E3 16 C3 FE
93 85 15 00 33 05 B8 00 13 86 F6 FF 63 54 D0 0C
33 07 A0 40 93 08 50 00 93 77 37 00 63 F4 C8 18
93 08 05 00 63 88 07 02 13 06 00 02 23 00 C5 00
13 77 27 00 63 00 07 14 13 07 F5 FF A3 00 C5 00
13 77 37 00 63 1A 07 14 23 01 C5 00 93 08 35 00
13 86 C6 FF 33 83 F6 40 B3 87 B7 00 B3 05 F8 00
13 77 C3 FF B7 27 20 20 33 07 B7 00 93 87 07 02
23 A0 F5 00 93 85 45 00 E3 9C E5 FE 93 77 33 00
63 88 07 04 13 73 C3 FF B3 87 68 00 33 06 66 40
13 07 00 02 23 80 E7 00 63 5C C0 02 A3 80 E7 00
93 05 10 00 63 06 B6 02 23 81 E7 00 93 05 20 00
63 00 B6 02 A3 81 E7 00 93 05 30 00 63 0A B6 00
23 82 E7 00 93 05 40 00 63 04 B6 00 A3 82 E7 00
33 05 D5 00 03 24 C1 05 83 24 81 05 13 01 01 06
67 80 00 00 13 04 00 00 6F F0 5F BF 93 F7 E7 FF
93 84 02 00 13 F5 27 00 93 0F 00 02 93 F3 07 02
E3 02 05 FE 6F F0 9F BB B3 05 B0 40 93 86 F6 FF
13 04 D0 02 E3 96 03 BC 93 87 05 00 13 05 00 00
13 03 C1 00 B3 F8 C7 02 93 05 05 00 13 05 15 00
B3 0E A3 00 13 8E 07 00 B3 08 1F 01 83 C8 08 00
B3 D7 C7 02 A3 8F 1E FF E3 7E CE FC 6F F0 DF BB
93 86 F6 FF 13 04 B0 02 6F F0 5F B8 93 07 00 03
23 00 F8 00 93 07 80 07 A3 00 F8 00 13 08 28 00
6F F0 9F CA 93 08 15 00 13 86 E6 FF 6F F0 9F ED
93 07 00 03 23 00 F8 00 13 08 18 00 6F F0 DF C8
93 86 E6 FF 6F F0 1F B6 93 08 25 00 13 86 D6 FF
6F F0 5F EB 93 07 05 00 6F F0 9F EE 93 07 08 00
6F F0 DF DE 93 86 0E 00 6F F0 1F C4 93 86 08 00
6F F0 1F D4 93 07 08 00 6F F0 5F CF 93 07 08 00
6F F0 1F BE
@4000174C
93 86 C1 1E 03 A7 06 00 B3 07 A7 00 23 A0 F6 00
13 85 01 1F 93 06 00 40 33 05 E5 00 63 D4 F6 00
73 00 10 00 67 80 00 00
@40001774
93 07 05 00 6F 00 80 01 03 C7 05 00 93 87 17 00
93 85 15 00 A3 8F E7 FE 63 04 07 08 33 E7 B7 00
13 77 37 00 E3 12 07 FE 83 A6 05 00 B7 08 FF FE
93 88 F8 EF 33 87 16 01 13 C6 F6 FF 37 88 80 80
33 77 C7 00 13 08 08 08 33 77 07 01 63 14 07 02
23 A0 D7 00 83 A6 45 00 93 87 47 00 93 85 45 00
33 87 16 01 13 C6 F6 FF 33 77 C7 00 33 77 07 01
E3 00 07 FE 23 80 D7 00 13 F7 F6 0F 63 02 07 02
13 D7 86 00 A3 80 E7 00 13 77 F7 0F 63 0A 07 00
13 D7 06 01 23 81 E7 00 13 77 F7 0F 63 14 07 00
67 80 00 00 93 D6 86 01 A3 81 D7 00 67 80 00 00
@40001824
B7 07 00 30 03 A5 07 00 67 80 00 00
@40001830
B7 07 00 20 03 A5 47 00 13 75 15 00 67 80 00 00
@40001840
37 07 00 20 83 27 47 00 93 F7 17 00 E3 9C 07 FE
93 07 A0 00 63 08 F5 00 B7 07 00 20 23 A6 A7 00
67 80 00 00 37 07 00 20 83 27 47 00 93 F7 17 00
E3 9C 07 FE 93 07 D0 00 23 26 F7 00 B7 07 00 20
23 A6 A7 00 67 80 00 00
@40001888
37 07 00 20 83 27 47 00 93 F7 17 00 E3 9C 07 FE
93 07 A0 00 63 08 F5 00 B7 07 00 20 23 A6 A7 00
67 80 00 00 37 07 00 20 83 27 47 00 93 F7 17 00
E3 9C 07 FE 93 07 D0 00 23 26 F7 00 B7 07 00 20
23 A6 A7 00 67 80 00 00
@400018D0
13 01 01 B7 23 20 21 47 23 26 11 46 23 24 81 46
23 22 91 46 23 2E 31 45 23 2C 41 45 23 2A 51 45
23 28 61 45 23 26 71 45 23 24 81 45 23 22 91 45
23 20 A1 45 23 2E B1 43 23 2A B1 46 23 2C C1 46
23 2E D1 46 23 20 E1 48 23 22 F1 48 23 24 01 49
23 26 11 49 83 47 05 00 13 09 41 47 23 2A 21 01
63 94 07 00 6F 10 00 09 13 0A 01 03 13 03 05 00
93 09 50 02 13 05 0A 00 93 04 00 01 13 84 C1 E3
13 0C 90 00 93 0B E0 02 13 0B C0 04 93 0A 70 03
63 82 37 0D 23 00 F5 00 83 47 13 00 13 05 15 00
13 03 13 00 E3 96 07 FE 23 00 05 00 83 46 01 03
63 94 06 00 6F 10 80 03 13 06 0A 00 37 07 00 20
93 05 A0 00 13 05 D0 00 83 27 47 00 93 F7 17 00
E3 9C 07 FE 63 8E B6 00 23 26 D7 00 83 46 16 00
93 07 16 00 63 86 06 02 13 86 07 00 6F F0 DF FD
83 27 47 00 93 F7 17 00 E3 9C 07 FE 23 26 A7 00
23 26 D7 00 83 46 16 00 93 07 16 00 E3 9E 06 FC
33 06 46 41 13 05 16 00 83 20 C1 46 03 24 81 46
83 24 41 46 03 29 01 46 83 29 C1 45 03 2A 81 45
83 2A 41 45 03 2B 01 45 83 2B C1 44 03 2C 81 44
83 2C 41 44 03 2D 01 44 83 2D C1 43 13 01 01 49
67 80 00 00 93 07 00 00 83 45 13 00 13 06 13 00
13 87 05 FE 13 77 F7 0F 63 EC E4 00 13 17 27 00
33 07 87 00 03 27 07 00 33 07 87 00 67 00 07 00
13 87 05 FD 13 77 F7 0F 63 78 EC 10 13 07 A0 02
93 06 F0 FF 63 8C E5 12 13 07 F0 FF 63 88 75 0D
13 F8 F5 0D 63 0C 68 09 13 88 F5 FB 13 78 F8 0F
63 EC 0A 05 93 88 01 E8 13 18 28 00 33 08 18 01
03 28 08 00 33 08 18 01 67 00 08 00 93 E7 17 00
13 03 06 00 6F F0 5F F8 93 E7 07 01 13 03 06 00
6F F0 9F F7 93 E7 47 00 13 03 06 00 6F F0 DF F6
93 E7 07 02 13 03 06 00 6F F0 1F F6 93 E7 87 00
13 03 06 00 6F F0 5F F5 93 0C 06 00 93 07 50 02
63 8A F5 00 23 00 F5 00 83 C5 0C 00 13 05 15 00
E3 84 05 E8 23 00 B5 00 83 C7 1C 00 13 83 1C 00
13 05 15 00 E3 9E 07 E4 6F F0 1F E7 93 88 05 00
83 45 16 00 93 0C 16 00 13 88 F5 FB 13 78 F8 0F
E3 EE 0A FB 13 83 01 F6 13 18 28 00 33 08 68 00
03 28 08 00 33 08 68 00 67 00 08 00 83 45 16 00
93 08 90 00 13 08 16 00 13 87 05 FD 13 77 F7 0F
63 F0 E8 7C 13 07 A0 02 63 8A E5 7E 13 06 08 00
13 07 00 00 6F F0 DF F0 93 06 00 00 13 08 90 00
13 97 26 00 33 07 D7 00 13 06 16 00 13 17 17 00
33 07 B7 00 83 45 06 00 93 06 07 FD 13 87 05 FD
13 77 F7 0F E3 7E E8 FC 6F F0 1F ED 83 26 09 00
83 45 23 00 13 06 23 00 13 09 49 00 E3 DE 06 EA
B3 06 D0 40 93 E7 07 01 6F F0 1F EB 93 E7 07 04
13 07 C0 06 63 84 E8 7A 83 28 09 00 13 09 49 00
03 C7 08 00 E3 1C 07 2A 13 07 00 03 93 05 10 00
23 0C E1 00 13 88 05 42 13 03 01 01 03 C7 18 00
33 03 68 00 13 08 E0 02 23 04 03 BF 13 06 20 00
E3 08 07 30 13 08 30 06 E3 50 E8 70 13 0E 40 06
33 6F C7 03 93 0E A0 00 13 06 06 42 93 0F 01 01
B3 0F F6 01 13 86 35 00 17 28 00 00 13 08 88 CD
33 47 C7 03 B3 45 DF 03 33 07 E8 00 03 47 07 00
23 84 EF BE 33 07 B8 00 83 45 07 00 33 67 DF 03
23 05 B3 BE 33 07 E8 00 03 48 07 00 93 05 01 01
13 07 06 42 B3 05 B7 00 13 07 16 00 23 84 05 BF
03 C6 28 00 93 05 07 42 13 08 01 01 33 83 05 01
93 05 E0 02 23 04 B3 BE 93 05 17 00 E3 0E 06 2A
13 08 30 06 E3 5C C8 62 13 0E 40 06 93 85 05 42
93 0F 01 01 B3 8F F5 01 93 05 37 00 93 0E A0 00
17 28 00 00 13 08 08 C5 33 6F C6 03 33 47 C6 03
33 46 DF 03 33 07 E8 00 03 47 07 00 23 84 EF BE
33 07 C8 00 33 66 DF 03 03 47 07 00 23 05 E3 BE
33 06 C8 00 03 48 06 00 13 87 05 42 13 06 01 01
33 06 C7 00 13 87 15 00 23 04 06 BF 93 05 07 42
03 C6 38 00 13 08 01 01 B3 88 05 01 93 05 E0 02
23 84 B8 BE 93 05 17 00 E3 04 06 26 13 08 30 06
E3 58 C8 56 13 03 40 06 93 85 05 42 13 0F 01 01
33 8F E5 01 93 05 37 00 13 0E A0 00 17 28 00 00
13 08 48 BC B3 6E 66 02 33 47 66 02 33 C6 CE 03
33 07 E8 00 03 47 07 00 23 04 EF BE 33 07 C8 00
33 E6 CE 03 03 47 07 00 23 85 E8 BE 33 06 C8 00
03 48 06 00 13 87 05 42 13 06 01 01 33 06 C7 00
23 04 06 BF 13 87 15 00 93 F7 07 01 63 9C 07 0C
13 88 F6 FF E3 5C D7 72 33 83 E6 40 B3 05 A0 40
93 08 F3 FF 13 06 50 00 93 F7 35 00 E3 78 16 73
13 06 05 00 63 88 07 02 13 08 00 02 23 00 05 01
93 F5 25 00 E3 8E 05 68 13 06 F5 FF A3 00 05 01
13 76 36 00 E3 18 06 60 23 01 05 01 13 06 35 00
13 88 C6 FF B3 08 F3 40 93 F5 C8 FF B3 07 F5 00
B7 26 20 20 B3 85 F5 00 93 86 06 02 23 A0 D7 00
93 87 47 00 E3 9C F5 FE 93 F6 C8 FF 93 F8 38 00
B3 07 D6 00 33 08 D8 40 63 82 08 04 93 06 00 02
23 80 D7 00 13 06 F8 FF 63 5A 07 03 A3 80 D7 00
93 05 E8 FF 63 54 C7 02 23 81 D7 00 13 06 D8 FF
63 5E B7 00 A3 81 D7 00 13 08 C8 FF 63 58 C7 00
23 82 D7 00 63 54 07 01 A3 82 D7 00 33 05 65 00
93 06 F7 FF 93 77 35 00 E3 84 07 36 83 47 E1 01
03 4E 81 01 03 43 91 01 83 48 A1 01 03 48 B1 01
83 45 C1 01 03 46 D1 01 23 03 F5 00 23 00 C5 01
A3 00 65 00 23 01 15 01 A3 01 05 01 23 02 B5 00
A3 02 C5 00 93 07 70 00 63 0E F7 06 03 46 F1 01
93 07 80 00 A3 03 C5 00 63 06 F7 06 03 46 01 02
93 07 90 00 23 04 C5 00 63 0E F7 04 03 46 11 02
93 07 A0 00 A3 04 C5 00 63 06 F7 04 03 46 21 02
93 07 B0 00 23 05 C5 00 63 0E F7 02 03 46 31 02
93 07 C0 00 A3 05 C5 00 63 06 F7 02 03 46 41 02
93 07 D0 00 23 06 C5 00 63 0E F7 00 03 46 51 02
93 07 F0 00 A3 06 C5 00 63 16 F7 00 83 47 61 02
23 07 F5 00 B3 08 E5 00 13 83 F6 FF E3 50 D7 52
33 88 E6 40 33 06 10 41 13 0E F8 FF 93 05 50 00
93 77 36 00 63 F8 C5 07 63 88 07 02 93 05 00 02
23 80 B8 00 13 76 26 00 E3 06 06 3E 13 86 F8 FF
A3 80 B8 00 13 76 36 00 E3 16 06 4C 23 81 B8 00
13 83 C6 FF 93 88 38 00 33 08 F8 40 B3 87 E7 00
B3 07 F5 00 93 75 C8 FF 37 26 20 20 B3 85 F5 00
13 06 06 02 23 A0 C7 00 93 87 47 00 E3 9C B7 FE
93 77 C8 FF 13 78 38 00 B3 88 F8 00 33 03 F3 40
63 02 08 04 13 06 00 02 23 80 C8 00 93 05 F3 FF
63 5A 67 02 A3 80 C8 00 93 07 E3 FF 63 54 B7 02
23 81 C8 00 93 05 D3 FF 63 5E F7 00 A3 81 C8 00
93 07 C3 FF 63 58 B7 00 23 82 C8 00 63 54 F7 00
A3 82 C8 00 33 05 D5 00 6F 00 C0 01 93 E7 07 04
13 06 00 01 13 08 49 00 83 25 09 00 13 09 08 00
EF F0 8F 9D 83 C7 1C 00 13 83 1C 00 E3 92 07 94
6F F0 9F 95 93 0C 06 00 93 F7 07 01 13 08 49 00
13 83 1C 00 63 8A 07 76 83 27 09 00 13 8E F6 FF
93 08 15 00 23 00 F5 00 E3 50 C0 51 33 07 10 41
13 86 E6 FF 93 0E 50 00 93 05 0E 00 93 77 37 00
63 D6 CE 06 63 86 07 02 13 0E 00 02 A3 00 C5 01
13 77 27 00 E3 0A 07 3A 23 01 C5 01 13 77 35 00
E3 10 07 3C A3 01 C5 01 93 08 45 00 13 8E C6 FF
B3 85 F5 40 93 87 17 00 B3 07 F5 00 13 F6 C5 FF
37 27 20 20 33 06 F6 00 13 07 07 02 23 A0 E7 00
93 87 47 00 E3 9C C7 FE 93 F7 C5 FF 93 F5 35 00
B3 88 F8 00 33 0E FE 40 63 84 05 04 93 07 00 02
23 80 F8 00 13 07 10 00 63 5C C7 03 A3 80 F8 00
13 07 20 00 63 06 EE 02 23 81 F8 00 13 07 30 00
63 00 EE 02 A3 81 F8 00 13 07 40 00 63 0A EE 00
23 82 F8 00 13 07 50 00 63 04 EE 00 A3 82 F8 00
83 C7 1C 00 33 05 D5 00 13 09 08 00 E3 92 07 84
6F F0 9F 85 93 0C 06 00 83 25 09 00 13 09 49 00
63 86 05 76 03 C6 05 00 E3 0E 06 24 E3 0C 07 24
13 86 05 00 6F 00 C0 00 33 08 E6 40 63 08 B8 00
03 48 16 00 13 06 16 00 E3 18 08 FE 93 F7 07 01
33 06 B6 40 63 82 07 74 63 56 C0 08 93 07 F6 FF
13 07 60 00 E3 70 F7 02 B3 E7 A5 00 93 F7 37 00
E3 9A 07 00 93 87 15 00 33 07 F5 40 13 37 37 00
E3 14 07 00 93 78 C6 FF 93 87 05 00 13 07 05 00
B3 88 B8 00 03 A8 07 00 93 87 47 00 13 07 47 00
23 2E 07 FF E3 98 F8 FE 93 77 C6 FF B3 85 F5 00
33 07 F5 00 63 06 F6 02 83 C8 05 00 13 88 17 00
23 00 17 01 63 5E C8 00 03 C8 15 00 93 87 27 00
A3 00 07 01 63 D6 C7 00 83 C7 25 00 23 01 F7 00
33 05 C5 00 13 8E F6 FF 13 83 1C 00 E3 50 D6 2C
B3 88 C6 40 33 07 A0 40 13 88 F8 FF 93 05 50 00
93 77 37 00 E3 F8 05 2D 13 08 05 00 63 80 07 04
93 05 00 02 23 00 B5 00 13 77 27 00 13 08 15 00
13 8E E6 FF 63 04 07 02 13 07 F5 FF A3 00 B5 00
13 77 37 00 13 08 25 00 13 8E D6 FF 63 18 07 00
13 08 35 00 23 01 B5 00 13 8E C6 FF B3 85 F8 40
93 F6 C5 FF B3 07 F5 00 37 27 20 20 B3 86 F6 00
13 07 07 02 23 A0 E7 00 93 87 47 00 E3 9C D7 FE
13 F7 C5 FF 93 F5 35 00 B3 07 E8 00 33 0E EE 40
63 82 05 04 93 06 00 02 23 80 D7 00 93 05 FE FF
63 5A C6 03 A3 80 D7 00 13 07 EE FF 63 54 B6 02
23 81 D7 00 93 05 DE FF 63 5E E6 00 A3 81 D7 00
13 07 CE FF 63 58 B6 00 23 82 D7 00 63 54 E6 00
A3 82 D7 00 83 C7 1C 00 33 05 15 01 63 92 07 E8
6F F0 8F E9 93 0C 06 00 13 06 F0 FF 63 88 C6 4A
83 25 09 00 13 06 00 01 13 09 49 00 EF E0 DF EE
83 C7 1C 00 13 83 1C 00 63 9C 07 E4 6F F0 CF E6
13 07 00 00 13 03 07 00 13 17 23 00 33 07 67 00
13 08 18 00 13 17 17 00 33 07 B7 00 83 45 08 00
13 03 07 FD 13 86 05 FD 13 76 F6 0F E3 FE C8 FC
13 07 03 00 13 06 08 00 6F F0 8F F2 03 27 09 00
83 45 26 00 13 09 49 00 13 48 F7 FF 13 58 F8 41
33 77 07 01 13 06 26 00 6F F0 8F F0 93 F5 07 04
17 17 00 00 13 07 07 59 63 86 05 00 17 17 00 00
13 07 C7 5A 03 28 09 00 93 05 A0 03 23 0D B1 00
83 48 08 00 83 43 18 00 83 4F 28 00 83 4E 38 00
03 43 48 00 13 FE F8 00 03 48 58 00 33 0E C7 01
93 D8 48 00 83 4D 0E 00 B3 08 17 01 93 DC 43 00
93 D2 4F 00 13 DF 4E 00 13 5E 43 00 93 F3 F3 00
93 FF FF 00 93 FE FE 00 13 73 F3 00 03 CD 08 00
B3 0C 97 01 B3 03 77 00 B3 02 57 00 B3 0F F7 01
33 0F E7 01 B3 0E D7 01 33 0E C7 01 33 03 67 00
93 58 48 00 83 CC 0C 00 83 C3 03 00 83 C2 02 00
83 CF 0F 00 03 4F 0F 00 83 CE 0E 00 03 4E 0E 00
03 43 03 00 B3 08 17 01 83 C8 08 00 93 9D 8D 00
33 6D BD 01 13 78 F8 00 23 1C A1 01 A3 0D 91 01
23 0E 71 00 A3 0E B1 00 23 0F 51 00 A3 0F F1 01
23 00 B1 02 A3 00 E1 03 23 01 D1 03 A3 01 B1 02
23 02 C1 03 A3 02 61 02 23 03 B1 02 33 07 07 01
A3 03 11 03 03 47 07 00 93 F7 07 01 23 26 E1 00
63 90 07 0E 93 07 10 01 93 85 F6 FF E3 D4 D7 0A
33 08 A0 40 13 87 E6 FE 93 0D 50 00 13 8D F6 FE
93 77 38 00 E3 F4 ED 08 13 07 05 00 63 88 07 02
93 05 00 02 23 00 B5 00 13 78 28 00 E3 08 08 02
13 07 F5 FF A3 00 B5 00 13 77 37 00 E3 1C 07 02
23 01 B5 00 13 07 35 00 93 85 C6 FF B3 0D FD 40
13 F8 CD FF B3 07 F5 00 B7 26 20 20 33 08 F8 00
93 86 06 02 23 A0 D7 00 93 87 47 00 E3 1C F8 FE
93 F7 CD FF 93 FD 3D 00 33 07 F7 00 B3 85 F5 40
63 84 0D 04 93 07 00 02 23 00 F7 00 93 06 10 01
63 DC B6 02 A3 00 F7 00 93 06 20 01 63 86 D5 02
23 01 F7 00 93 06 30 01 63 80 D5 02 A3 01 F7 00
93 06 40 01 63 8A D5 00 23 02 F7 00 93 06 50 01
63 84 D5 00 A3 02 F7 00 33 05 A5 01 93 06 00 01
93 77 35 00 63 94 07 70 83 27 C1 01 23 22 F5 00
83 27 01 02 23 24 F5 00 83 27 81 01 23 20 F5 00
83 27 41 02 23 26 F5 00 83 27 C1 00 13 08 15 01
93 88 F6 FF 23 08 F5 00 93 07 10 01 63 DC D7 72
33 07 00 41 93 85 E6 FE 13 0E 50 00 13 83 F6 FE
93 77 37 00 63 7E BE 06 63 8E 07 02 93 05 00 02
A3 08 B5 00 13 77 27 00 13 08 25 01 93 88 E6 FF
63 02 07 02 23 09 B5 00 13 77 35 00 13 08 35 01
93 88 D6 FF 63 18 07 00 13 08 45 01 A3 09 B5 00
93 88 C6 FF 33 03 F3 40 93 87 17 01 B3 07 F5 00
93 75 C3 FF 37 27 20 20 B3 85 F5 00 13 07 07 02
23 A0 E7 00 93 87 47 00 E3 9C B7 FE 93 77 C3 FF
13 73 33 00 33 08 F8 00 B3 88 F8 40 63 04 03 04
93 07 00 02 23 00 F8 00 13 07 10 01 63 5C 17 03
A3 00 F8 00 13 07 20 01 63 86 E8 02 23 01 F8 00
13 07 30 01 63 80 E8 02 A3 01 F8 00 13 07 40 01
63 8A E8 00 23 02 F8 00 13 07 50 01 63 84 E8 00
A3 02 F8 00 33 05 D5 00 83 47 26 00 13 09 49 00
13 03 26 00 63 9E 07 AC 6F F0 0F AF 13 06 30 06
63 54 E6 3C 13 03 40 06 B3 6F 67 02 13 0F A0 00
17 18 00 00 13 08 08 26 13 06 40 00 93 05 30 00
13 0E 20 00 B3 CE EF 03 33 47 67 02 33 03 D8 01
83 4E 03 00 93 9E 8E 00 33 07 E8 00 03 43 07 00
33 E7 EF 03 33 63 D3 01 23 1C 61 00 33 07 E8 00
03 47 07 00 13 08 0E 42 13 03 01 01 33 0E 68 00
23 04 EE BE 13 88 05 42 13 03 01 01 03 C7 18 00
33 03 68 00 13 08 E0 02 23 04 03 BF 63 1C 07 CE
13 07 06 42 13 06 01 01 33 06 C7 00 13 87 25 00
93 05 00 03 23 04 B6 BE 13 08 01 01 93 05 07 42
03 C6 28 00 33 83 05 01 93 05 E0 02 23 04 B3 BE
93 05 17 00 63 16 06 D4 13 86 05 42 93 05 01 01
33 06 B6 00 13 07 27 00 93 05 00 03 23 04 B6 BE
13 08 01 01 93 05 07 42 03 C6 38 00 B3 88 05 01
93 05 E0 02 23 84 B8 BE 93 05 17 00 63 10 06 DA
13 86 05 42 93 05 01 01 33 06 B6 00 93 05 00 03
13 07 27 00 23 04 B6 BE 6F F0 0F DF 93 E7 17 00
93 06 80 00 6F F0 DF B4 93 07 10 00 63 DE D7 44
13 86 F6 FF B3 05 A0 40 93 88 E6 FF 13 07 50 00
93 0E 06 00 93 F7 35 00 63 5A 17 55 13 07 05 00
63 88 07 02 13 06 00 02 23 00 C5 00 93 F5 25 00
63 8C 05 50 13 07 F5 FF A3 00 C5 00 13 77 37 00
63 10 07 52 23 01 C5 00 13 07 35 00 13 86 C6 FF
B3 85 FE 40 13 FE C5 FF B3 07 F5 00 B7 28 20 20
33 0E FE 00 93 88 08 02 23 A0 17 01 93 87 47 00
E3 1C FE FE 93 F8 C5 FF 93 F5 35 00 B3 07 17 01
33 06 16 41 63 84 05 04 13 07 00 02 23 80 E7 00
93 05 10 00 63 DC C5 02 A3 80 E7 00 93 05 20 00
63 06 B6 02 23 81 E7 00 93 05 30 00 63 00 B6 02
A3 81 E7 00 93 05 40 00 63 0A B6 00 23 82 E7 00
93 05 50 00 63 04 B6 00 A3 82 E7 00 83 27 09 00
B3 0E D5 01 33 05 D5 00 23 80 FE 00 83 C7 1C 00
13 09 08 00 63 96 07 8C 6F F0 0F 8E 97 15 00 00
93 85 45 0B 6F F0 9F 89 13 87 F6 FF 63 5A D6 34
33 8E C6 40 B3 08 A0 40 13 03 FE FF 13 08 50 00
93 F7 38 00 63 70 68 46 13 08 05 00 63 8C 07 02
13 03 00 02 23 00 65 00 93 F8 28 00 13 08 15 00
13 87 E6 FF 63 80 08 02 13 07 F5 FF A3 00 65 00
13 77 37 00 63 14 07 44 13 08 35 00 23 01 65 00
13 87 C6 FF B3 06 FE 40 13 F3 C6 FF B3 07 F5 00
B7 28 20 20 33 03 F3 00 93 88 08 02 23 A0 17 01
93 87 47 00 E3 1C F3 FE 93 F8 C6 FF 93 F6 36 00
B3 07 18 01 33 07 17 41 63 82 06 04 93 06 00 02
23 80 D7 00 13 08 F7 FF 63 5A E6 02 A3 80 D7 00
93 08 E7 FF 63 54 06 03 23 81 D7 00 13 08 D7 FF
63 5E 16 01 A3 81 D7 00 13 07 C7 FF 63 58 06 01
23 82 D7 00 63 54 E6 00 A3 82 D7 00 33 05 C5 01
93 06 F6 FF 6F F0 4F FE 93 E7 27 00 13 06 A0 00
6F F0 4F E7 93 87 15 00 B3 85 C5 00 13 07 05 00
6F 00 80 00 93 87 17 00 03 C8 F7 FF 13 07 17 00
A3 0F 07 FF E3 98 B7 FE 6F F0 9F 83 13 05 00 00
6F F0 8F 82 13 0A 01 03 13 05 0A 00 6F E0 DF FA
83 25 81 01 93 57 27 00 13 06 10 00 23 20 B5 00
63 8A C7 26 83 25 C1 01 13 06 30 00 23 22 B5 00
63 96 C7 00 83 27 01 02 23 24 F5 00 93 77 37 00
63 82 07 D2 93 77 C7 FF 33 06 F5 00 13 08 01 01
93 85 07 42 B3 85 05 01 03 C8 85 BE 93 85 17 00
23 00 06 01 63 D0 E5 D0 93 85 17 42 13 08 01 01
B3 85 05 01 83 C5 85 BE 93 87 27 00 A3 00 B6 00
63 D2 E7 CE 93 87 07 42 B3 87 07 01 83 C7 87 BE
23 01 F6 00 6F F0 0F CD 13 06 90 00 63 54 E6 10
93 0E A0 00 33 43 D7 03 17 18 00 00 13 08 88 E9
13 06 30 00 93 05 20 00 13 0E 10 00 33 03 68 00
03 43 03 00 33 67 D7 03 23 0C 61 00 6F F0 1F C5
93 08 90 00 17 18 00 00 13 08 C8 E6 63 D8 C8 AC
13 03 A0 00 B3 48 66 02 93 85 05 42 13 0E 01 01
33 8E C5 01 93 05 27 00 33 07 18 01 03 47 07 00
33 66 66 02 23 04 EE BE 6F F0 4F AA 13 03 90 00
17 18 00 00 13 08 08 E3 63 54 C3 A0 13 0E A0 00
33 43 C6 03 93 85 05 42 93 0E 01 01 B3 8E D5 01
93 05 27 00 33 07 68 00 03 47 07 00 33 66 C6 03
23 84 EE BE 6F F0 CF 9D 13 03 90 00 17 18 00 00
13 08 48 DF 63 50 E3 94 13 0E A0 00 33 43 C7 03
13 06 06 42 93 0E 01 01 B3 0E D6 01 13 86 25 00
B3 05 68 00 83 C5 05 00 33 67 C7 03 23 84 BE BE
6F F0 4F 91 93 88 18 00 13 83 E6 FF 6F F0 CF C2
93 0C 06 00 93 E7 27 00 13 08 49 00 13 06 A0 00
6F F0 8F CA 13 06 20 00 93 05 10 00 13 0E 00 00
17 18 00 00 13 08 08 D9 6F F0 5F B6 13 06 80 00
6F F0 4F C8 13 06 A0 00 6F F0 CF C7 93 0C 06 00
6F F0 8F 83 13 F6 07 01 E3 08 06 D0 13 06 00 00
6F F0 4F E5 93 0C 06 00 13 08 49 00 13 06 80 00
6F F0 8F C5 93 0C 06 00 93 E7 07 04 13 08 49 00
13 06 00 01 6F F0 4F C4 93 0C 06 00 13 08 49 00
13 06 00 01 6F F0 4F C3 93 E7 07 04 93 0C 06 00
6F E0 9F FE 13 06 25 00 13 88 D6 FF 6F F0 8F 9F
93 0C 06 00 13 08 49 00 13 06 A0 00 6F F0 CF C0
93 06 07 00 6F F0 4F D6 83 27 09 00 13 05 15 00
13 09 08 00 A3 0F F5 FE 83 C7 1C 00 63 84 07 00
6F E0 1F D4 6F E0 5F D5 93 08 25 00 13 0E 06 00
6F F0 0F C6 93 88 28 00 13 83 D6 FF 6F F0 CF B3
93 08 35 00 13 8E D6 FF 6F F0 8F C4 13 85 08 00
6F F0 4F BC 13 06 45 00 93 07 40 00 6F F0 1F DB
13 06 15 00 13 88 E6 FF 6F F0 CF 97 83 45 81 01
03 47 91 01 93 07 A0 03 23 00 B5 00 A3 00 E5 00
23 01 F5 00 A3 01 95 01 23 02 75 00 A3 02 F5 00
23 03 55 00 A3 03 F5 01 23 04 F5 00 A3 04 E5 01
23 05 D5 01 A3 05 F5 00 23 06 C5 01 A3 06 65 00
23 07 F5 00 A3 07 15 01 6F F0 1F 8D 83 C7 1C 00
63 84 07 00 6F E0 DF C9 6F E0 1F CB 93 06 08 00
6F F0 4F 99 13 05 08 00 6F F0 1F 9A 93 07 05 00
6F F0 CF 93 93 07 05 00 6F F0 CF DA 13 07 15 00
93 85 E6 FF 6F F0 8F FE 13 07 15 00 13 86 08 00
6F F0 1F B0 13 07 25 00 93 85 D6 FF 6F F0 0F FD
13 07 25 00 13 86 D6 FF 6F F0 9F AE 93 07 05 00
6F F0 9F B1 93 07 05 00 6F F0 5F C1 13 07 05 00
6F F0 4F FE 93 86 05 00 6F F0 9F 82 13 08 25 00
13 87 D6 FF 6F F0 1F BC 13 85 08 00 6F F0 1F B4
@40002D50
B7 07 08 02 93 87 17 00 37 07 00 20 23 20 F7 00
67 80 00 00
@40002D64
B7 07 00 30 83 A7 07 00 23 A4 F1 1E 67 80 00 00
@40002D74
B7 07 00 30 83 A7 07 00 23 A2 F1 1E 67 80 00 00
@40002D84
03 A5 41 1E 83 A7 81 1E 33 05 F5 40 67 80 00 00
@40002D94
13 01 01 FF 23 26 11 00 EF D0 1F BA 97 17 00 00
93 87 07 B5 03 A6 07 00 83 A6 47 00 EF D0 8F CC
83 20 C1 00 13 01 01 01 67 80 00 00
@40002DC0
13 01 01 FF 23 20 21 01 13 89 01 1E 83 27 09 00
23 24 81 00 03 24 05 00 83 A6 07 00 03 AF 47 00
83 AE 87 00 03 AE 07 01 03 A3 47 01 83 A8 87 01
03 A8 C7 01 83 A5 47 02 03 A6 87 02 03 A7 C7 02
23 26 11 00 23 22 91 00 93 04 05 00 03 A5 07 02
23 20 D4 00 83 A6 04 00 23 22 E4 01 23 24 D4 01
23 28 C4 01 23 2A 64 00 23 2C 14 01 23 2E 04 01
23 20 A4 02 23 22 B4 02 23 24 C4 02 23 26 E4 02
13 07 50 00 23 A6 E4 00 23 20 D4 00 83 A7 07 00
23 26 E4 00 83 A5 81 1D 23 20 F4 00 03 26 09 00
13 05 A0 00 13 06 C6 00 EF 00 10 19 83 27 44 00
63 80 07 08 83 A7 04 00 83 20 C1 00 03 24 81 00
83 AF 07 00 03 AF 47 00 83 AE 87 00 03 AE C7 00
03 A3 07 01 83 A8 47 01 03 A8 87 01 83 A5 C7 01
03 A6 07 02 83 A6 47 02 03 A7 87 02 83 A7 C7 02
23 A0 F4 01 23 A2 E4 01 23 A4 D4 01 23 A6 C4 01
23 A8 64 00 23 AA 14 01 23 AC 04 01 23 AE B4 00
23 A0 C4 02 23 A2 D4 02 23 A4 E4 02 23 A6 F4 02
03 29 01 00 83 24 41 00 13 01 01 01 67 80 00 00
03 A5 84 00 93 07 60 00 93 05 84 00 23 26 F4 00
EF 00 90 0A 83 27 09 00 03 25 C4 00 13 06 C4 00
83 A7 07 00 83 20 C1 00 83 24 41 00 23 20 F4 00
03 24 81 00 03 29 01 00 93 05 A0 00 13 01 01 01
6F 00 90 0C
@40002F34
13 01 01 F6 B7 07 08 02 93 87 17 00 37 07 00 20
23 2E 11 08 23 2C 81 08 23 2A 91 08 23 28 21 09
23 26 31 09 23 24 41 09 23 22 51 09 23 20 61 09
23 2E 71 07 23 2C 81 07 23 2A 91 07 23 28 A1 07
23 26 B1 07 23 20 F7 00 17 15 00 00 13 05 C5 A1
EF E0 DF 94 13 87 C1 1E 83 27 07 00 93 86 01 1F
93 05 00 40 13 86 07 03 23 20 C7 00 B3 86 F6 00
63 D4 C5 00 73 00 10 00 83 27 07 00 13 8D C1 1D
23 20 DD 00 93 86 07 03 23 20 D7 00 13 86 01 1F
13 07 00 40 B3 07 F6 00 63 54 D7 00 73 00 10 00
03 27 0D 00 13 85 07 01 23 A2 07 00 23 A0 E7 00
13 07 20 00 23 A4 E7 00 13 07 80 02 23 A6 E7 00
97 15 00 00 93 85 85 9B 93 8C 01 1E 23 A0 FC 00
EF E0 0F F7 97 15 00 00 93 85 45 9C 13 05 01 02
EF E0 0F F6 93 07 A0 00 17 17 00 00 13 07 C7 78
17 15 00 00 13 05 45 BD 23 2E F7 64 EF E0 1F 8A
17 15 00 00 13 05 85 9B EF E0 5F 89 17 15 00 00
13 05 85 BB EF E0 9F 88 83 A7 C1 1C 63 8A 07 6A
17 15 00 00 13 05 85 9C EF E0 5F 87 17 15 00 00
13 05 85 B9 EF E0 9F 86 B7 85 1E 00 93 85 05 48
17 15 00 00 13 05 45 A0 B7 5A 52 59 B7 04 FF FE
37 84 80 80 EF E0 9F 84 93 09 10 00 13 8B 11 1D
93 8B 41 1D 13 89 01 1D 13 8C 81 1D 93 8A 4A 84
93 84 F4 EF 13 04 04 08 93 07 10 04 23 00 FB 00
93 07 10 00 23 A0 FB 00 93 07 20 04 23 00 F9 00
93 06 01 04 13 87 0A 00 17 16 00 00 13 06 C6 88
13 06 46 00 23 A0 E6 00 03 27 06 00 93 86 46 00
B3 07 97 00 93 45 F7 FF B3 F7 B7 00 B3 F7 87 00
E3 80 07 FE 23 80 E6 00 93 77 F7 0F 63 86 07 02
93 57 87 00 A3 80 F6 00 93 F7 F7 0F 63 8E 07 00
93 57 07 01 23 81 F6 00 93 F7 F7 0F 63 86 07 00
13 57 87 01 A3 81 E6 00 93 07 10 00 93 05 01 04
13 05 01 02 23 2E F1 00 EF 00 00 75 93 37 15 00
13 06 81 01 93 05 30 00 23 A0 FB 00 13 05 20 00
93 07 70 00 23 2C F1 00 EF 00 C0 69 83 26 81 01
13 06 30 00 97 15 00 00 93 85 05 64 13 85 01 5F
EF 00 40 69 03 A5 0C 00 EF F0 5F C4 03 47 09 00
93 07 00 04 63 F6 E7 54 93 0D 10 04 13 0A 30 00
6F 00 40 01 03 47 09 00 93 87 1D 00 93 FD F7 0F
63 62 B7 0B 93 05 30 04 13 85 0D 00 EF 00 C0 6B
03 27 C1 01 E3 10 E5 FE 93 05 C1 01 13 05 00 00
EF 00 40 5E 13 06 01 04 93 86 0A 00 97 05 00 00
93 85 85 7A 93 85 45 00 23 20 D6 00 83 A6 05 00
13 06 46 00 33 87 96 00 13 C5 F6 FF 33 77 A7 00
33 77 87 00 E3 00 07 FE 23 00 D6 00 13 F7 F6 0F
63 06 07 02 13 D7 86 00 A3 00 E6 00 13 77 F7 0F
63 0E 07 00 13 D7 06 01 23 01 E6 00 13 77 F7 0F
63 06 07 00 93 D6 86 01 A3 01 D6 00 03 47 09 00
93 87 1D 00 23 20 3C 01 93 FD F7 0F 13 8A 09 00
E3 72 B7 F7 93 17 1A 00 33 8A 47 01 03 28 81 01
83 46 0B 00 93 07 10 04 33 46 0A 03 13 07 06 00
63 98 F6 00 83 27 0C 00 13 07 96 00 33 07 F7 40
B7 87 1E 00 93 89 19 00 93 87 17 48 E3 96 F9 E2
B7 07 00 30 83 A7 07 00 03 A4 81 1E 17 15 00 00
13 05 85 81 33 84 87 40 23 26 E1 00 23 24 C1 00
23 22 01 01 23 A2 F1 1E 23 A2 81 1C EF E0 0F E2
17 15 00 00 13 05 45 94 EF E0 4F E1 17 05 00 00
13 05 85 7F EF E0 8F E0 17 15 00 00 13 05 C5 92
EF E0 CF DF 83 25 0C 00 17 15 00 00 13 05 45 81
EF E0 CF DE 93 05 50 00 17 15 00 00 13 05 05 82
EF E0 CF DD 83 A5 0B 00 17 15 00 00 13 05 C5 82
EF E0 CF DC 93 05 10 00 17 15 00 00 13 05 05 80
EF E0 CF DB 83 45 0B 00 17 15 00 00 13 05 85 82
EF E0 CF DA 93 05 10 04 17 15 00 00 13 05 45 83
EF E0 CF D9 83 45 09 00 17 15 00 00 13 05 05 84
EF E0 CF D8 93 05 20 04 17 15 00 00 13 05 45 81
EF E0 CF D7 93 87 01 1F 83 A5 07 42 17 15 00 00
13 05 85 83 EF E0 8F D6 93 05 70 00 17 05 00 00
13 05 C5 79 EF E0 8F D5 97 17 00 00 93 87 C7 42
83 A5 C7 65 17 15 00 00 13 05 C5 82 EF E0 0F D4
17 15 00 00 13 05 C5 83 EF E0 4F D3 17 15 00 00
13 05 C5 85 EF E0 8F D2 83 A7 0C 00 17 15 00 00
13 05 85 85 83 A5 07 00 EF E0 4F D1 17 15 00 00
13 05 45 86 EF E0 8F D0 83 A7 0C 00 17 15 00 00
13 05 85 88 83 A5 47 00 EF E0 4F CF 93 05 00 00
17 05 00 00 13 05 85 72 EF E0 4F CE 83 A7 0C 00
17 15 00 00 13 05 05 88 83 A5 87 00 EF E0 0F CD
93 05 20 00 17 05 00 00 13 05 45 70 EF E0 0F CC
83 A7 0C 00 17 15 00 00 13 05 85 87 83 A5 C7 00
EF E0 CF CA 93 05 10 01 17 05 00 00 13 05 05 6E
EF E0 CF C9 83 A5 0C 00 17 15 00 00 13 05 05 87
93 85 05 01 EF E0 8F C8 17 15 00 00 13 05 C5 87
EF E0 CF C7 17 15 00 00 13 05 85 8A EF E0 0F C7
83 27 0D 00 17 05 00 00 13 05 05 7A 83 A5 07 00
EF E0 CF C5 17 15 00 00 13 05 C5 89 EF E0 0F C5
83 27 0D 00 17 05 00 00 13 05 05 7D 83 A5 47 00
EF E0 CF C3 93 05 00 00 17 05 00 00 13 05 05 67
EF E0 CF C2 83 27 0D 00 17 05 00 00 13 05 85 7C
83 A5 87 00 EF E0 8F C1 93 05 10 00 17 05 00 00
13 05 C5 64 EF E0 8F C0 83 27 0D 00 17 05 00 00
13 05 05 7C 83 A5 C7 00 EF E0 4F BF 93 05 20 01
17 05 00 00 13 05 85 62 EF E0 4F BE 83 25 0D 00
17 05 00 00 13 05 85 7B 93 85 05 01 EF E0 0F BD
17 05 00 00 13 05 45 7C EF E0 4F BC 03 27 C1 00
17 15 00 00 13 05 05 84 93 05 07 00 EF E0 0F BB
93 05 50 00 17 05 00 00 13 05 45 5E EF E0 0F BA
03 28 41 00 03 26 81 00 17 15 00 00 13 05 45 83
33 0A 0A 41 93 15 3A 00 B3 85 45 41 B3 85 C5 40
EF E0 CF B7 93 05 D0 00 17 05 00 00 13 05 05 5B
EF E0 CF B6 83 25 81 01 17 15 00 00 13 05 05 82
EF E0 CF B5 93 05 70 00 17 05 00 00 13 05 05 59
EF E0 CF B4 83 25 C1 01 17 15 00 00 13 05 C5 81
EF E0 CF B3 93 05 10 00 17 05 00 00 13 05 05 57
EF E0 CF B2 93 05 01 02 17 15 00 00 13 05 85 81
EF E0 CF B1 17 15 00 00 13 05 85 82 EF E0 0F B1
93 05 01 04 17 15 00 00 13 05 05 85 EF E0 0F B0
17 15 00 00 13 05 05 86 EF E0 4F AF 17 05 00 00
13 05 85 61 EF E0 8F AE 23 A0 81 1C 93 07 10 00
63 D4 87 0E 13 05 04 00 EF D0 1F A9 97 05 00 00
83 A5 85 2F 13 04 05 00 EF D0 CF ED 97 05 00 00
83 A5 C5 2E EF D0 4F BA 93 07 05 00 93 84 C1 1B
93 05 04 00 17 05 00 00 03 25 45 2D 23 A0 F4 00
EF D0 8F B8 93 07 05 00 13 84 81 1B 17 15 00 00
13 05 45 88 23 20 F4 00 EF E0 4F A8 03 A5 04 00
EF D0 9F 9C 93 05 05 00 17 15 00 00 13 05 85 89
EF E0 CF A6 17 15 00 00 13 05 45 89 EF E0 0F A6
03 25 04 00 EF D0 5F 9A 93 05 05 00 17 15 00 00
13 05 45 87 EF E0 8F A4 17 05 00 00 13 05 C5 56
EF E0 CF A3 83 20 C1 09 03 24 81 09 83 24 41 09
03 29 01 09 83 29 C1 08 03 2A 81 08 83 2A 41 08
03 2B 01 08 83 2B C1 07 03 2C 81 07 83 2C 41 07
03 2D 01 07 83 2D C1 06 13 01 01 0A 67 80 00 00
13 0A 90 00 6F F0 9F B7 17 05 00 00 13 05 05 79
EF E0 CF 9E 17 05 00 00 13 05 C5 7B EF E0 0F 9E
17 05 00 00 13 05 45 50 EF E0 4F 9D 6F F0 9F F9
17 05 00 00 13 05 45 34 EF E0 4F 9C 17 05 00 00
13 05 85 4E EF E0 8F 9B 6F F0 1F 95
@40003720
03 C7 11 1D 93 07 10 04 63 04 F7 00 67 80 00 00
83 27 05 00 03 A7 81 1D 93 87 97 00 B3 87 E7 40
23 20 F5 00 67 80 00 00
@40003748
93 87 01 1E 03 A6 07 00 63 08 06 00 03 27 06 00
23 20 E5 00 03 A6 07 00 13 06 C6 00 83 A5 81 1D
13 05 A0 00 6F 00 C0 08
@40003770
13 87 41 1D 83 26 07 00 83 C7 11 1D 93 87 F7 FB
93 B7 17 00 B3 E7 D7 00 23 20 F7 00 93 07 20 04
23 88 F1 1C 67 80 00 00
@40003798
93 07 10 04 A3 88 F1 1C 23 AA 01 1C 67 80 00 00
@400037A8
93 07 20 00 63 00 F5 04 13 07 30 00 23 A0 E5 00
13 07 10 00 63 0A E5 00 13 07 40 00 63 00 E5 02
63 0A 05 00 67 80 00 00 03 A7 81 1D 93 07 40 06
E3 DA E7 FE 23 A0 05 00 67 80 00 00 23 A0 F5 00
67 80 00 00 93 07 10 00 23 A0 F5 00 67 80 00 00
@400037F8
13 05 25 00 B3 05 B5 00 23 20 B6 00 67 80 00 00
@40003808
13 07 56 00 13 08 80 0C 33 08 07 03 13 16 26 00
93 17 27 00 33 05 F5 00 23 20 D5 00 23 2C E5 06
23 22 D5 00 B3 07 C8 00 B3 87 F5 00 83 A6 07 01
23 AA E7 00 23 AC E7 00 13 87 16 00 23 A8 E7 00
03 27 05 00 B3 85 05 01 B3 85 C5 00 B7 17 00 00
B3 87 B7 00 23 AA E7 FA 93 07 50 00 23 AC F1 1C
67 80 00 00
@4000386C
13 75 F5 0F 93 F5 F5 0F 63 06 B5 00 13 05 00 00
67 80 00 00 A3 88 A1 1C 13 05 10 00 67 80 00 00
@4000388C
13 01 01 FF 23 26 11 00 83 47 25 00 03 C7 35 00
13 06 00 00 93 06 00 00 63 8A E7 02 63 84 06 00
A3 88 C1 1C EF C0 DF 84 93 07 00 00 63 58 A0 00
93 07 A0 00 23 AC F1 1C 93 07 10 00 83 20 C1 00
13 85 07 00 13 01 01 01 67 80 00 00 93 06 10 00
13 86 07 00 6F F0 5F FC
@400038E4
13 05 E5 FF 13 35 15 00 67 80 00 00
@400038F0
00 00 00 00 38 9C 8C 41 00 24 74 49 5B 47 DA 56
@40003900
30 31 32 33 34 35 36 37 38 39 61 62 63 64 65 66
67 68 69 6A 6B 6C 6D 6E 6F 70 71 72 73 74 75 76
77 78 79 7A 00 00 00 00 30 31 32 33 34 35 36 37
38 39 41 42 43 44 45 46 47 48 49 4A 4B 4C 4D 4E
4F 50 51 52 53 54 55 56 57 58 59 5A 00 00 00 00
3C 4E 55 4C 4C 3E 00 00 44 48 52 59 53 54 4F 4E
45 20 50 52 4F 47 52 41 4D 2C 20 32 27 4E 44 20
53 54 52 49 4E 47 00 00 44 48 52 59 53 54 4F 4E
45 20 50 52 4F 47 52 41 4D 2C 20 33 27 52 44 20
53 54 52 49 4E 47 00 00 44 68 72 79 73 74 6F 6E
65 20 42 65 6E 63 68 6D 61 72 6B 00 44 48 52 59
53 54 4F 4E 45 20 50 52 4F 47 52 41 4D 2C 20 53
4F 4D 45 20 53 54 52 49 4E 47 00 00 44 48 52 59
53 54 4F 4E 45 20 50 52 4F 47 52 41 4D 2C 20 31
27 53 54 20 53 54 52 49 4E 47 00 00 44 68 72 79
73 74 6F 6E 65 20 42 65 6E 63 68 6D 61 72 6B 2C
20 56 65 72 73 69 6F 6E 20 32 2E 31 20 28 4C 61
6E 67 75 61 67 65 3A 20 43 29 0A 00 50 72 6F 67
72 61 6D 20 63 6F 6D 70 69 6C 65 64 20 77 69 74
68 20 27 72 65 67 69 73 74 65 72 27 20 61 74 74
72 69 62 75 74 65 0A 00 50 72 6F 67 72 61 6D 20
63 6F 6D 70 69 6C 65 64 20 77 69 74 68 6F 75 74
20 27 72 65 67 69 73 74 65 72 27 20 61 74 74 72
69 62 75 74 65 0A 00 00 45 78 65 63 75 74 69 6F
6E 20 73 74 61 72 74 73 2C 20 25 64 20 72 75 6E
73 20 74 68 72 6F 75 67 68 20 44 68 72 79 73 74
6F 6E 65 0A 00 00 00 00 45 78 65 63 75 74 69 6F
6E 20 65 6E 64 73 0A 00 46 69 6E 61 6C 20 76 61
6C 75 65 73 20 6F 66 20 74 68 65 20 76 61 72 69
61 62 6C 65 73 20 75 73 65 64 20 69 6E 20 74 68
65 20 62 65 6E 63 68 6D 61 72 6B 3A 0A 00 00 00
49 6E 74 5F 47 6C 6F 62 3A 20 20 20 20 20 20 20
20 20 20 20 20 25 64 0A 00 00 00 00 20 20 20 20
20 20 20 20 73 68 6F 75 6C 64 20 62 65 3A 20 20
20 25 64 0A 00 00 00 00 42 6F 6F 6C 5F 47 6C 6F
62 3A 20 20 20 20 20 20 20 20 20 20 20 25 64 0A
00 00 00 00 43 68 5F 31 5F 47 6C 6F 62 3A 20 20
20 20 20 20 20 20 20 20 20 25 63 0A 00 00 00 00
20 20 20 20 20 20 20 20 73 68 6F 75 6C 64 20 62
65 3A 20 20 20 25 63 0A 00 00 00 00 43 68 5F 32
5F 47 6C 6F 62 3A 20 20 20 20 20 20 20 20 20 20
20 25 63 0A 00 00 00 00 41 72 72 5F 31 5F 47 6C
6F 62 5B 38 5D 3A 20 20 20 20 20 20 20 25 64 0A
00 00 00 00 41 72 72 5F 32 5F 47 6C 6F 62 5B 38
5D 5B 37 5D 3A 20 20 20 20 25 64 0A 00 00 00 00
20 20 20 20 20 20 20 20 73 68 6F 75 6C 64 20 62
65 3A 20 20 20 4E 75 6D 62 65 72 5F 4F 66 5F 52
75 6E 73 20 2B 20 31 30 0A 00 00 00 50 74 72 5F
47 6C 6F 62 2D 3E 0A 00 20 20 50 74 72 5F 43 6F
6D 70 3A 20 20 20 20 20 20 20 20 20 20 25 64 0A
00 00 00 00 20 20 20 20 20 20 20 20 73 68 6F 75
6C 64 20 62 65 3A 20 20 20 28 69 6D 70 6C 65 6D
65 6E 74 61 74 69 6F 6E 2D 64 65 70 65 6E 64 65
6E 74 29 0A 00 00 00 00 20 20 44 69 73 63 72 3A
20 20 20 20 20 20 20 20 20 20 20 20 20 25 64 0A
00 00 00 00 20 20 45 6E 75 6D 5F 43 6F 6D 70 3A
20 20 20 20 20 20 20 20 20 25 64 0A 00 00 00 00
20 20 49 6E 74 5F 43 6F 6D 70 3A 20 20 20 20 20
20 20 20 20 20 25 64 0A 00 00 00 00 20 20 53 74
72 5F 43 6F 6D 70 3A 20 20 20 20 20 20 20 20 20
20 25 73 0A 00 00 00 00 20 20 20 20 20 20 20 20
73 68 6F 75 6C 64 20 62 65 3A 20 20 20 44 48 52
59 53 54 4F 4E 45 20 50 52 4F 47 52 41 4D 2C 20
53 4F 4D 45 20 53 54 52 49 4E 47 0A 00 00 00 00
4E 65 78 74 5F 50 74 72 5F 47 6C 6F 62 2D 3E 0A
00 00 00 00 20 20 20 20 20 20 20 20 73 68 6F 75
6C 64 20 62 65 3A 20 20 20 28 69 6D 70 6C 65 6D
65 6E 74 61 74 69 6F 6E 2D 64 65 70 65 6E 64 65
6E 74 29 2C 20 73 61 6D 65 20 61 73 20 61 62 6F
76 65 0A 00 49 6E 74 5F 31 5F 4C 6F 63 3A 20 20
20 20 20 20 20 20 20 20 20 25 64 0A 00 00 00 00
49 6E 74 5F 32 5F 4C 6F 63 3A 20 20 20 20 20 20
20 20 20 20 20 25 64 0A 00 00 00 00 49 6E 74 5F
33 5F 4C 6F 63 3A 20 20 20 20 20 20 20 20 20 20
20 25 64 0A 00 00 00 00 45 6E 75 6D 5F 4C 6F 63
3A 20 20 20 20 20 20 20 20 20 20 20 20 25 64 0A
00 00 00 00 53 74 72 5F 31 5F 4C 6F 63 3A 20 20
20 20 20 20 20 20 20 20 20 25 73 0A 00 00 00 00
20 20 20 20 20 20 20 20 73 68 6F 75 6C 64 20 62
65 3A 20 20 20 44 48 52 59 53 54 4F 4E 45 20 50
52 4F 47 52 41 4D 2C 20 31 27 53 54 20 53 54 52
49 4E 47 0A 00 00 00 00 53 74 72 5F 32 5F 4C 6F
63 3A 20 20 20 20 20 20 20 20 20 20 20 25 73 0A
00 00 00 00 20 20 20 20 20 20 20 20 73 68 6F 75
6C 64 20 62 65 3A 20 20 20 44 48 52 59 53 54 4F
4E 45 20 50 52 4F 47 52 41 4D 2C 20 32 27 4E 44
20 53 54 52 49 4E 47 0A 00 00 00 00 4D 65 61 73
75 72 65 64 20 74 69 6D 65 20 74 6F 6F 20 73 6D
61 6C 6C 20 74 6F 20 6F 62 74 61 69 6E 20 6D 65
61 6E 69 6E 67 66 75 6C 20 72 65 73 75 6C 74 73
0A 00 00 00 50 6C 65 61 73 65 20 69 6E 63 72 65
61 73 65 20 6E 75 6D 62 65 72 20 6F 66 20 72 75
6E 73 0A 00 4D 69 63 72 6F 73 65 63 6F 6E 64 73
20 66 6F 72 20 6F 6E 65 20 72 75 6E 20 74 68 72
6F 75 67 68 20 44 68 72 79 73 74 6F 6E 65 3A 20
00 00 00 00 25 64 20 0A 00 00 00 00 44 68 72 79
73 74 6F 6E 65 73 20 70 65 72 20 53 65 63 6F 6E
64 3A 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 00
@40003F2C
A0 DB FF FF 24 DB FF FF 24 DB FF FF 94 DB FF FF
24 DB FF FF 24 DB FF FF 24 DB FF FF 24 DB FF FF
24 DB FF FF 24 DB FF FF 24 DB FF FF 88 DB FF FF
24 DB FF FF 7C DB FF FF 24 DB FF FF 24 DB FF FF
70 DB FF FF 68 EC FF FF 68 DB FF FF 68 DB FF FF
68 DB FF FF 68 DB FF FF 68 DB FF FF 68 DB FF FF
68 DB FF FF 68 DB FF FF 68 DB FF FF 68 DB FF FF
68 DB FF FF 68 DB FF FF 68 DB FF FF 68 DB FF FF
68 DB FF FF 68 DB FF FF 68 DB FF FF 68 DB FF FF
68 DB FF FF 68 DB FF FF 68 DB FF FF 68 DB FF FF
44 EC FF FF 68 DB FF FF 68 DB FF FF 68 DB FF FF
68 DB FF FF 68 DB FF FF 68 DB FF FF 68 DB FF FF
68 DB FF FF 1C EC FF FF 68 DB FF FF B4 E0 FF FF
E0 EB FF FF 68 DB FF FF 68 DB FF FF 68 DB FF FF
68 DB FF FF E0 EB FF FF 68 DB FF FF 68 DB FF FF
68 DB FF FF 68 DB FF FF 68 DB FF FF 34 EC FF FF
74 E3 FF FF 68 DB FF FF 68 DB FF FF B4 E1 FF FF
68 DB FF FF 80 EC FF FF 68 DB FF FF 68 DB FF FF
58 EC FF FF 6C DB FF FF 8C DA FF FF 8C DA FF FF
8C DA FF FF 8C DA FF FF 8C DA FF FF 8C DA FF FF
8C DA FF FF 8C DA FF FF 8C DA FF FF 8C DA FF FF
8C DA FF FF 8C DA FF FF 8C DA FF FF 8C DA FF FF
8C DA FF FF 8C DA FF FF 8C DA FF FF 8C DA FF FF
8C DA FF FF 8C DA FF FF 8C DA FF FF 8C DA FF FF
AC DF FF FF 8C DA FF FF 8C DA FF FF 8C DA FF FF
8C DA FF FF 8C DA FF FF 8C DA FF FF 8C DA FF FF
8C DA FF FF 70 DB FF FF 8C DA FF FF D8 DF FF FF
38 E9 FF FF 8C DA FF FF 8C DA FF FF 8C DA FF FF
8C DA FF FF 38 E9 FF FF 8C DA FF FF 8C DA FF FF
8C DA FF FF 8C DA FF FF 8C DA FF FF 2C EB FF FF
98 E2 FF FF 8C DA FF FF 8C DA FF FF D8 E0 FF FF
8C DA FF FF 34 EB FF FF 8C DA FF FF 8C DA FF FF
B0 DF FF FF 1C 09 00 40 CC 04 00 40 44 08 00 40
CC 04 00 40 08 09 00 40 CC 04 00 40 44 08 00 40
1C 09 00 40 1C 09 00 40 08 09 00 40 44 08 00 40
A8 04 00 40 A8 04 00 40 A8 04 00 40 08 09 00 40
DC 0C 00 40 1C 0B 00 40 60 0C 00 40 1C 0B 00 40
CC 0C 00 40 1C 0B 00 40 60 0C 00 40 DC 0C 00 40
DC 0C 00 40 CC 0C 00 40 60 0C 00 40 F8 0A 00 40
F8 0A 00 40 F8 0A 00 40 CC 0C 00 40 00 01 02 02
03 03 03 03 04 04 04 04 04 04 04 04 05 05 05 05
05 05 05 05 05 05 05 05 05 05 05 05 06 06 06 06
06 06 06 06 06 06 06 06 06 06 06 06 06 06 06 06
06 06 06 06 06 06 06 06 06 06 06 06 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08
