// MIKROISLEM KODLARININ PARCALARI
// MI[7]...MI[0] Ilgili birime girecek mi girmeyecek mi onu gosteriyor
// Onundeki 5 bit ise o birime giren hangi buyruk oldugunu belirtiyor
// Simdilik toplam 15 bit

// MI[0]
`define AMBVAR 1'b1
`define AMBYOK 1'b0

// MI[1]
`define CLAVAR 1'b1
`define CLAYOK 1'b0

// MI[2]
`define BDCVAR 1'b1
`define BDCYOK 1'b0

// MI[3]
`define BIBVAR 1'b1
`define BIBYOK 1'b0

// MI[4]
`define DALVAR 1'b1
`define DALYOK 1'b0

// MI[5]
`define SIFVAR 1'b1
`define SIFYOK 1'b0

// MI[6]
`define YAPVAR 1'b1
`define YAPYOK 1'b0

// MI[7]
`define SISVAR 1'b1
`define SISYOK 1'b0

// IMM ve CMP ilk 5 bitin icine yedirilebilir, bit sayisi azalir
// Cozden sonraki asamalarda compressed olmasinin onemi kalmayacaksa burada tamamen kaldirabiliriz, bu nasil cozdugumuze bagli

// MI[8]
`define IMMVAR 1'b1
`define IMMYOK 1'b0

// MI[9]
`define CMPVAR 1'b1
`define CMPYOK 1'b0

// MIKROISLEM KODLARI
// Toplam 87 buyruk

`define GECERSIZ 15'b00000_00_00000000

// AMB buyruklari
`define AND_MI   {5'b0_0_0_0_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define AUIPC_MI {5'b0_0_0_0_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR} 
`define LUI_MI   {5'b0_0_0_1_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}  
`define OR_MI    {5'b0_0_0_1_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR} 
`define SLL_MI   {5'b0_0_1_0_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}  
`define SLT_MI   {5'b0_0_1_0_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}  
`define SLTU_MI  {5'b0_0_1_1_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}   
`define SRA_MI   {5'b0_0_1_1_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}  
`define SRL_MI   {5'b0_1_0_0_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}  
`define XOR_MI   {5'b0_1_0_0_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}  

// IMMLI AMB buyruklari
`define ANDI_MI  {5'b0_1_0_1_0, CMPYOK, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define ORI_MI   {5'b0_1_0_1_1, CMPYOK, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define SLLI_MI  {5'b0_1_1_0_0, CMPYOK, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define SLTI_MI  {5'b0_1_1_0_1, CMPYOK, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define SLTIU_MI {5'b0_1_1_1_0, CMPYOK, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define SRAI_MI  {5'b0_1_1_1_1, CMPYOK, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define SRLI_MI  {5'b1_0_0_0_0, CMPYOK, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define XORI_MI  {5'b1_0_0_0_1, CMPYOK, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}

// Compressed AMB buyruklari
`define C_AND_MI {5'b1_0_0_1_0, CMPVAR, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define C_OR_MI  {5'b1_0_0_1_1, CMPVAR, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define C_XOR_MI {5'b1_0_1_0_0, CMPVAR, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}

// Compressed IMMLI AMB buyruklari
`define C_ANDI_MI {5'b1_0_1_0_0, CMPVAR, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define C_SLLI_MI {5'b1_0_1_0_1, CMPVAR, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define C_SRAI_MI {5'b1_0_1_1_0, CMPVAR, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define C_SRLI_MI {5'b1_0_1_1_1, CMPVAR, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}

// Bolme buyruklari, simdilik amb'de olsun?
`define DIV_MI  {5'b1_1_0_0_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define DIVU_MI {5'b1_1_0_0_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define REM_MI  {5'b1_1_0_1_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}
`define REMU_MI {5'b1_1_0_1_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBVAR}

// Carry Lookahead Toplayici buyruklari
`define ADD_MI {5'b0_0_0_0_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAVAR, AMBYOK}
`define SUB_MI {5'b0_0_0_0_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAVAR, AMBYOK}
// cikarmayi amb'ye mi almaliyiz?

// Carry Lookahead IMMLI Toplayici buyruklari
`define ADDI_MI {5'b0_0_0_1_0, CMPYOK, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAVAR, AMBYOK}

// Compressed Carry Lookahead Toplayici buyruklari
`define C_ADD_MI {5'b0_0_0_1_1, CMPVAR, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAVAR, AMBYOK}
`define C_MV_MI  {5'b0_0_1_0_0, CMPVAR, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAVAR, AMBYOK}
`define C_SUB_MI {5'b0_0_1_0_1, CMPVAR, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAVAR, AMBYOK}

// Compressed IMMLI Carry Lookahead Toplayici buyruklari
`define C_ADDI_MI     {5'b0_0_1_1_0, CMPVAR, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAVAR, AMBYOK}
`define C_ADDI16SP_MI {5'b0_0_1_1_1, CMPVAR, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAVAR, AMBYOK}
`define C_ADDI4SPN_MI {5'b0_1_0_0_0, CMPVAR, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAVAR, AMBYOK}
`define C_LI_MI       {5'b0_1_0_0_1, CMPVAR, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAVAR, AMBYOK}
`define C_NOP_MI      {5'b0_1_0_1_0, CMPVAR, IMMVAR, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAVAR, AMBYOK}

// Modified Booth Dadda Carpici buyruklari
`define MUL_MI    {5'b0_0_0_0_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCVAR, CLAYOK, AMBYOK}
`define MULH_MI   {5'b0_0_0_0_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCVAR, CLAYOK, AMBYOK}
`define MULHSU_MI {5'b0_0_0_1_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCVAR, CLAYOK, AMBYOK}
`define MULHU_MI  {5'b0_0_0_1_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCVAR, CLAYOK, AMBYOK}

// BIB buyruklari
`define LB_MI  {5'b0_0_0_0_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}
`define LBU_MI {5'b0_0_0_0_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}
`define LH_MI  {5'b0_0_0_1_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}
`define LHU_MI {5'b0_0_0_1_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}
`define LW_MI  {5'b0_0_1_0_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}

`define SB_MI  {5'b0_0_1_0_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}
`define SH_MI  {5'b0_0_1_1_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}
`define SW_MI  {5'b0_0_1_1_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}

// Compressed BIB buyruklari
`define C_LUI_MI  {5'b0_1_0_0_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}
`define C_LW_MI   {5'b0_1_0_0_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}
`define C_LWSP_MI {5'b0_1_0_1_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}
`define C_SW_MI   {5'b0_1_0_1_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}
`define C_SWSP_MI {5'b0_1_1_0_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}

// Out-of-order BIB buyruklari
// Bizim islemci in-order oldugu icin bu buyruklari implement etmemize gerek yok, bos birakin
`define FENCE_MI   {5'b0_1_1_0_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}
`define FENCE_I_MI {5'b0_1_1_1_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALYOK, BIBVAR, BDCYOK, CLAYOK, AMBYOK}

// Dallanma buyruklari
`define BEQ_MI  {5'b0_0_0_0_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALVAR, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define BGE_MI  {5'b0_0_0_0_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALVAR, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define BGEU_MI {5'b0_0_0_1_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALVAR, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define BLT_MI  {5'b0_0_0_1_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALVAR, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define BLTU_MI {5'b0_0_1_0_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALVAR, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define BNE_MI  {5'b0_0_1_0_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALVAR, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define JAL_MI  {5'b0_0_1_1_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALVAR, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define JALR_MI {5'b0_0_1_1_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALVAR, BIBYOK, BDCYOK, CLAYOK, AMBYOK}

// Compressed Dallanma buyruklari
`define C_BEQZ_MI {5'b0_1_0_0_0, CMPVAR, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALVAR, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define C_BNEZ_MI {5'b0_1_0_0_1, CMPVAR, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALVAR, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define C_J_MI    {5'b0_1_0_1_0, CMPVAR, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALVAR, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define C_JAL_MI  {5'b0_1_0_1_1, CMPVAR, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALVAR, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define C_JALR_MI {5'b0_1_1_0_0, CMPVAR, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALVAR, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define C_JR_MI   {5'b0_1_1_0_1, CMPVAR, IMMYOK, SISYOK, YAPYOK, SIFYOK, DALVAR, BIBYOK, BDCYOK, CLAYOK, AMBYOK}

// Sifreleme buyruklari
`define HMDST_MI {5'b0_0_0_0_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFVAR, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define PKG_MI   {5'b0_0_0_0_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFVAR, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define RVRS_MI  {5'b0_0_0_1_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFVAR, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define SLADD_MI {5'b0_0_0_1_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFVAR, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define CNTZ_MI  {5'b0_0_1_0_0, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFVAR, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define CNTP_MI  {5'b0_0_1_0_1, CMPYOK, IMMYOK, SISYOK, YAPYOK, SIFVAR, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBYOK}

// Yapay Zeka buyruklari
`define CONV_LD_W_MI  {5'b0_0_0_0_0, CMPYOK, IMMYOK, SISYOK, YAPVAR, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define CONV_CLR_W_MI {5'b0_0_0_0_1, CMPYOK, IMMYOK, SISYOK, YAPVAR, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define CONV_LD_X_MI  {5'b0_0_0_1_0, CMPYOK, IMMYOK, SISYOK, YAPVAR, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define CONV_CLR_X_MI {5'b0_0_0_1_1, CMPYOK, IMMYOK, SISYOK, YAPVAR, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define CONV_RUN_MI   {5'b0_0_1_0_0, CMPYOK, IMMYOK, SISYOK, YAPVAR, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBYOK}

// Sistem buyruklari
`define EBREAK_MI {5'b0_0_0_0_0, CMPYOK, IMMYOK, SISVAR, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
`define ECALL_MI  {5'b0_0_0_0_0, CMPYOK, IMMYOK, SISVAR, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBYOK}

// Compressed Sistem buyruklari
`define C_EBREAK_MI {5'b0_0_0_0_0, CMPVAR, IMMYOK, SISVAR, YAPYOK, SIFYOK, DALYOK, BIBYOK, BDCYOK, CLAYOK, AMBYOK}
