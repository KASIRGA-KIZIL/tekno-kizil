// zero_counter.v


`timescale 1ns / 1ps


module zero_counter(
    input [31:0] deger_i,
    output reg [4:0] sifir_sayisi,
    output [0:0] hepsi_sifir
);
    assign hepsi_sifir = !(|deger_i);
    always@*begin
        sifir_sayisi = 5'd0;
        casez(deger_i)
            32'b10000000_00000000_00000000_00000000:
                sifir_sayisi = 5'd31;
            32'b?1000000_00000000_00000000_00000000:
                sifir_sayisi = 5'd30;
            32'b??100000_00000000_00000000_00000000:
                sifir_sayisi = 5'd29;
            32'b???10000_00000000_00000000_00000000:
                sifir_sayisi = 5'd28;
            32'b????1000_00000000_00000000_00000000:
                sifir_sayisi = 5'd27;
            32'b?????100_00000000_00000000_00000000:
                sifir_sayisi = 5'd26;
            32'b??????10_00000000_00000000_00000000:
                sifir_sayisi = 5'd25;
            32'b???????1_00000000_00000000_00000000:
                sifir_sayisi = 5'd24;
            32'b????????_10000000_00000000_00000000:
                sifir_sayisi = 5'd23;
            32'b????????_?1000000_00000000_00000000:
                sifir_sayisi = 5'd22;
            32'b????????_??100000_00000000_00000000:
                sifir_sayisi = 5'd21;
            32'b????????_???10000_00000000_00000000:
                sifir_sayisi = 5'd20;
            32'b????????_????1000_00000000_00000000:
                sifir_sayisi = 5'd19;
            32'b????????_?????100_00000000_00000000:
                sifir_sayisi = 5'd18;
            32'b????????_??????10_00000000_00000000:
                sifir_sayisi = 5'd17;
            32'b????????_???????1_00000000_00000000:
                sifir_sayisi = 5'd16;
            32'b????????_????????_10000000_00000000:
                sifir_sayisi = 5'd15;
            32'b????????_????????_?1000000_00000000:
                sifir_sayisi = 5'd14;
            32'b????????_????????_??100000_00000000:
                sifir_sayisi = 5'd13;
            32'b????????_????????_???10000_00000000:
                sifir_sayisi = 5'd12;
            32'b????????_????????_????1000_00000000:
                sifir_sayisi = 5'd11;
            32'b????????_????????_?????100_00000000:
                sifir_sayisi = 5'd10;
            32'b????????_????????_??????10_00000000:
                sifir_sayisi = 5'd9;
            32'b????????_????????_???????1_00000000:
                sifir_sayisi = 5'd8;
            32'b????????_????????_????????_10000000:
                sifir_sayisi = 5'd7;
            32'b00000000_????????_????????_?1000000:
                sifir_sayisi = 5'd6;
            32'b????????_????????_????????_??100000:
                sifir_sayisi = 5'd5;
            32'b????????_????????_????????_???10000:
                sifir_sayisi = 5'd4;
            32'b????????_????????_????????_????1000:
                sifir_sayisi = 5'd3;
            32'b????????_????????_????????_?????100:
                sifir_sayisi = 5'd2;
            32'b????????_????????_????????_??????10:
                sifir_sayisi = 5'd1;
            32'b????????_????????_????????_???????1:
                sifir_sayisi = 5'd0;
        endcase
    end
endmodule
