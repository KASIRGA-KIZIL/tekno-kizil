// getir.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module getir(
    input clk_i,
    input rst_i


);


endmodule
