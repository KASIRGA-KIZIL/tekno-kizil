// veri_onbellegi_denetleyicisi.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module veri_onbellegi_denetleyicisi(
    input clk_i,
    input rst_i


);


endmodule
