// tb_bellek_islem_birimi.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module tb_bellek_islem_birimi();

    bellek_islem_birimi bib(

    );

    initial begin

        $finish;
    end

endmodule
