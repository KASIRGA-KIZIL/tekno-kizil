module progmem (
    // Closk & reset
    input wire clk,
    input wire rstn,

    // PicoRV32 bus interface
    input  wire        valid,
    output wire        ready,
    input  wire [31:0] addr,
    output wire [31:0] rdata
);

  // ============================================================================

  localparam MEM_SIZE_BITS = 10;  // In 32-bit words
  localparam MEM_SIZE = 1 << MEM_SIZE_BITS;
  localparam MEM_ADDR_MASK = 32'h0010_0000;

  // ============================================================================

  wire [MEM_SIZE_BITS-1:0] mem_addr;
  reg  [             31:0] mem_data;
  reg  [             31:0] mem      [0:MEM_SIZE];

  initial begin

  mem['h0000] <= 32'hff010113;
  mem['h0001] <= 32'h00112623;
  mem['h0002] <= 32'h00812423;
  mem['h0003] <= 32'h3c5000ef;
  mem['h0004] <= 32'h00001517;
  mem['h0005] <= 32'hc0450513;
  mem['h0006] <= 32'h2dc000ef;
  mem['h0007] <= 32'h00001517;
  mem['h0008] <= 32'hc0050513;
  mem['h0009] <= 32'h2d0000ef;
  mem['h000A] <= 32'h3d1000ef;
  mem['h000B] <= 32'h3cd000ef;
  mem['h000C] <= 32'h3c9000ef;
  mem['h000D] <= 32'h3c5000ef;
  mem['h000E] <= 32'h00001517;
  mem['h000F] <= 32'hbec50513;
  mem['h0010] <= 32'h2b4000ef;
  mem['h0011] <= 32'h00001417;
  mem['h0012] <= 32'hbe440413;
  mem['h0013] <= 32'h3ad000ef;
  mem['h0014] <= 32'h00050593;
  mem['h0015] <= 32'h00040513;
  mem['h0016] <= 32'h29c000ef;
  mem['h0017] <= 32'hff1ff06f;
  mem['h0018] <= 32'h0000006f;
  mem['h0019] <= 32'hfa010113;
  mem['h001A] <= 32'h04812e23;
  mem['h001B] <= 32'h04912c23;
  mem['h001C] <= 32'h0407f813;
  mem['h001D] <= 32'h00001e97;
  mem['h001E] <= 32'hbe0e8e93;
  mem['h001F] <= 32'h00081663;
  mem['h0020] <= 32'h00001e97;
  mem['h0021] <= 32'hbace8e93;
  mem['h0022] <= 32'h0107f413;
  mem['h0023] <= 32'h14041663;
  mem['h0024] <= 32'h0017f813;
  mem['h0025] <= 32'h0117f493;
  mem['h0026] <= 32'h03000393;
  mem['h0027] <= 32'h14080263;
  mem['h0028] <= 32'h0027f813;
  mem['h0029] <= 32'h0207ff13;
  mem['h002A] <= 32'h12080463;
  mem['h002B] <= 32'h1405c463;
  mem['h002C] <= 32'h0047f813;
  mem['h002D] <= 32'h18081463;
  mem['h002E] <= 32'h0087f793;
  mem['h002F] <= 32'h00000f93;
  mem['h0030] <= 32'h00078663;
  mem['h0031] <= 32'hfff68693;
  mem['h0032] <= 32'h02000f93;
  mem['h0033] <= 32'h000f0c63;
  mem['h0034] <= 32'h01000793;
  mem['h0035] <= 32'h18f60e63;
  mem['h0036] <= 32'hff860793;
  mem['h0037] <= 32'h0017b793;
  mem['h0038] <= 32'h40f686b3;
  mem['h0039] <= 32'h12059063;
  mem['h003A] <= 32'h03000793;
  mem['h003B] <= 32'h00f10623;
  mem['h003C] <= 32'h00100813;
  mem['h003D] <= 32'h00c10293;
  mem['h003E] <= 32'h00080893;
  mem['h003F] <= 32'h00e85463;
  mem['h0040] <= 32'h00070893;
  mem['h0041] <= 32'h411686b3;
  mem['h0042] <= 32'h02049063;
  mem['h0043] <= 32'h00d50733;
  mem['h0044] <= 32'h02000793;
  mem['h0045] <= 32'h16d05a63;
  mem['h0046] <= 32'h00150513;
  mem['h0047] <= 32'hfef50fa3;
  mem['h0048] <= 32'hfee51ce3;
  mem['h0049] <= 32'hfff00693;
  mem['h004A] <= 32'h000f8663;
  mem['h004B] <= 32'h01f50023;
  mem['h004C] <= 32'h00150513;
  mem['h004D] <= 32'h000f0a63;
  mem['h004E] <= 32'h00800793;
  mem['h004F] <= 32'h12f60263;
  mem['h0050] <= 32'h01000793;
  mem['h0051] <= 32'h10f60263;
  mem['h0052] <= 32'h00041e63;
  mem['h0053] <= 32'h00d507b3;
  mem['h0054] <= 32'h14d05063;
  mem['h0055] <= 32'h00150513;
  mem['h0056] <= 32'hfe750fa3;
  mem['h0057] <= 32'hfea79ce3;
  mem['h0058] <= 32'hfff00693;
  mem['h0059] <= 32'h410887b3;
  mem['h005A] <= 32'h00f507b3;
  mem['h005B] <= 32'h03000713;
  mem['h005C] <= 32'h11185863;
  mem['h005D] <= 32'h00150513;
  mem['h005E] <= 32'hfee50fa3;
  mem['h005F] <= 32'hfea79ce3;
  mem['h0060] <= 32'h00b28733;
  mem['h0061] <= 32'h00078613;
  mem['h0062] <= 32'h00074803;
  mem['h0063] <= 32'h00070513;
  mem['h0064] <= 32'h00160613;
  mem['h0065] <= 32'hff060fa3;
  mem['h0066] <= 32'hfff70713;
  mem['h0067] <= 32'hfea296e3;
  mem['h0068] <= 32'h00158593;
  mem['h0069] <= 32'h00b785b3;
  mem['h006A] <= 32'h0cd05863;
  mem['h006B] <= 32'h00d58533;
  mem['h006C] <= 32'h02000793;
  mem['h006D] <= 32'h00158593;
  mem['h006E] <= 32'hfef58fa3;
  mem['h006F] <= 32'hfeb51ce3;
  mem['h0070] <= 32'h05c12403;
  mem['h0071] <= 32'h05812483;
  mem['h0072] <= 32'h06010113;
  mem['h0073] <= 32'h00008067;
  mem['h0074] <= 32'h00000f93;
  mem['h0075] <= 32'hef9ff06f;
  mem['h0076] <= 32'hffe7f793;
  mem['h0077] <= 32'h00040493;
  mem['h0078] <= 32'h0027f813;
  mem['h0079] <= 32'h02000393;
  mem['h007A] <= 32'h0207ff13;
  mem['h007B] <= 32'hfe0802e3;
  mem['h007C] <= 32'hebdff06f;
  mem['h007D] <= 32'h40b005b3;
  mem['h007E] <= 32'hfff68693;
  mem['h007F] <= 32'h02d00f93;
  mem['h0080] <= 32'hec0f18e3;
  mem['h0081] <= 32'h00058793;
  mem['h0082] <= 32'h00000813;
  mem['h0083] <= 32'h00c10293;
  mem['h0084] <= 32'h02c7f8b3;
  mem['h0085] <= 32'h00080593;
  mem['h0086] <= 32'h00180813;
  mem['h0087] <= 32'h01028e33;
  mem['h0088] <= 32'h00078313;
  mem['h0089] <= 32'h011e88b3;
  mem['h008A] <= 32'h0008c883;
  mem['h008B] <= 32'h02c7d7b3;
  mem['h008C] <= 32'hff1e0fa3;
  mem['h008D] <= 32'hfcc37ee3;
  mem['h008E] <= 32'hec1ff06f;
  mem['h008F] <= 32'hfff68693;
  mem['h0090] <= 32'h02b00f93;
  mem['h0091] <= 32'he89ff06f;
  mem['h0092] <= 32'h03000793;
  mem['h0093] <= 32'h00f50023;
  mem['h0094] <= 32'h07800793;
  mem['h0095] <= 32'h00f500a3;
  mem['h0096] <= 32'h00250513;
  mem['h0097] <= 32'heedff06f;
  mem['h0098] <= 32'h03000793;
  mem['h0099] <= 32'h00f50023;
  mem['h009A] <= 32'h00150513;
  mem['h009B] <= 32'heddff06f;
  mem['h009C] <= 32'hffe68693;
  mem['h009D] <= 32'he71ff06f;
  mem['h009E] <= 32'h00058513;
  mem['h009F] <= 32'hf45ff06f;
  mem['h00A0] <= 32'h00050793;
  mem['h00A1] <= 32'hefdff06f;
  mem['h00A2] <= 32'hfff68693;
  mem['h00A3] <= 32'he9dff06f;
  mem['h00A4] <= 32'hfff68693;
  mem['h00A5] <= 32'hed1ff06f;
  mem['h00A6] <= 32'h20000737;
  mem['h00A7] <= 32'h00472783;
  mem['h00A8] <= 32'h0017f793;
  mem['h00A9] <= 32'hfe079ce3;
  mem['h00AA] <= 32'h00a70623;
  mem['h00AB] <= 32'h00008067;
  mem['h00AC] <= 32'h00054683;
  mem['h00AD] <= 32'h02068263;
  mem['h00AE] <= 32'h20000737;
  mem['h00AF] <= 32'h00150513;
  mem['h00B0] <= 32'h00472783;
  mem['h00B1] <= 32'h0017f793;
  mem['h00B2] <= 32'hfe079ce3;
  mem['h00B3] <= 32'h00d70623;
  mem['h00B4] <= 32'h00054683;
  mem['h00B5] <= 32'hfe0694e3;
  mem['h00B6] <= 32'h00008067;
  mem['h00B7] <= 32'h20000737;
  mem['h00B8] <= 32'h00472783;
  mem['h00B9] <= 32'h0017f793;
  mem['h00BA] <= 32'hfe079ce3;
  mem['h00BB] <= 32'h00a70623;
  mem['h00BC] <= 32'h00008067;
  mem['h00BD] <= 32'hb7010113;
  mem['h00BE] <= 32'h48e12023;
  mem['h00BF] <= 32'h46112623;
  mem['h00C0] <= 32'h46812423;
  mem['h00C1] <= 32'h46912223;
  mem['h00C2] <= 32'h47212023;
  mem['h00C3] <= 32'h45312e23;
  mem['h00C4] <= 32'h45412c23;
  mem['h00C5] <= 32'h45512a23;
  mem['h00C6] <= 32'h45612823;
  mem['h00C7] <= 32'h45712623;
  mem['h00C8] <= 32'h45812423;
  mem['h00C9] <= 32'h45912223;
  mem['h00CA] <= 32'h45a12023;
  mem['h00CB] <= 32'h43b12e23;
  mem['h00CC] <= 32'h46b12a23;
  mem['h00CD] <= 32'h46c12c23;
  mem['h00CE] <= 32'h46d12e23;
  mem['h00CF] <= 32'h48f12223;
  mem['h00D0] <= 32'h49012423;
  mem['h00D1] <= 32'h49112623;
  mem['h00D2] <= 32'h00054783;
  mem['h00D3] <= 32'h47410713;
  mem['h00D4] <= 32'h00e12a23;
  mem['h00D5] <= 32'h72078a63;
  mem['h00D6] <= 32'h03010993;
  mem['h00D7] <= 32'h00050313;
  mem['h00D8] <= 32'h00070a13;
  mem['h00D9] <= 32'h00098513;
  mem['h00DA] <= 32'h02500913;
  mem['h00DB] <= 32'h01000493;
  mem['h00DC] <= 32'h00001417;
  mem['h00DD] <= 32'h91440413;
  mem['h00DE] <= 32'h00900d93;
  mem['h00DF] <= 32'h02e00c93;
  mem['h00E0] <= 32'h04c00d13;
  mem['h00E1] <= 32'h03700c13;
  mem['h00E2] <= 32'h05278863;
  mem['h00E3] <= 32'h00f50023;
  mem['h00E4] <= 32'h00134783;
  mem['h00E5] <= 32'h00150513;
  mem['h00E6] <= 32'h00130313;
  mem['h00E7] <= 32'hfe0796e3;
  mem['h00E8] <= 32'h00050023;
  mem['h00E9] <= 32'h03014603;
  mem['h00EA] <= 32'h10060863;
  mem['h00EB] <= 32'h00098693;
  mem['h00EC] <= 32'h20000737;
  mem['h00ED] <= 32'h00472783;
  mem['h00EE] <= 32'h0017f793;
  mem['h00EF] <= 32'hfe079ce3;
  mem['h00F0] <= 32'h00c70623;
  mem['h00F1] <= 32'h0016c603;
  mem['h00F2] <= 32'h00168793;
  mem['h00F3] <= 32'h12060463;
  mem['h00F4] <= 32'h00078693;
  mem['h00F5] <= 32'hfe1ff06f;
  mem['h00F6] <= 32'h00000793;
  mem['h00F7] <= 32'h00134603;
  mem['h00F8] <= 32'h00130593;
  mem['h00F9] <= 32'hfe060713;
  mem['h00FA] <= 32'h0ff77713;
  mem['h00FB] <= 32'h00e4ec63;
  mem['h00FC] <= 32'h00271713;
  mem['h00FD] <= 32'h00870733;
  mem['h00FE] <= 32'h00072703;
  mem['h00FF] <= 32'h00870733;
  mem['h0100] <= 32'h00070067;
  mem['h0101] <= 32'hfd060713;
  mem['h0102] <= 32'h0ff77713;
  mem['h0103] <= 32'h14edfc63;
  mem['h0104] <= 32'h02a00713;
  mem['h0105] <= 32'hfff00693;
  mem['h0106] <= 32'h18e60063;
  mem['h0107] <= 32'hfff00713;
  mem['h0108] <= 32'h11960c63;
  mem['h0109] <= 32'h0df67813;
  mem['h010A] <= 32'h09a80c63;
  mem['h010B] <= 32'hfbf60813;
  mem['h010C] <= 32'h0ff87813;
  mem['h010D] <= 32'h050c6e63;
  mem['h010E] <= 32'h00001897;
  mem['h010F] <= 32'h89088893;
  mem['h0110] <= 32'h00281813;
  mem['h0111] <= 32'h01180833;
  mem['h0112] <= 32'h00082803;
  mem['h0113] <= 32'h01180833;
  mem['h0114] <= 32'h00080067;
  mem['h0115] <= 32'h0017e793;
  mem['h0116] <= 32'h00058313;
  mem['h0117] <= 32'hf81ff06f;
  mem['h0118] <= 32'h0107e793;
  mem['h0119] <= 32'h00058313;
  mem['h011A] <= 32'hf75ff06f;
  mem['h011B] <= 32'h0047e793;
  mem['h011C] <= 32'h00058313;
  mem['h011D] <= 32'hf69ff06f;
  mem['h011E] <= 32'h0207e793;
  mem['h011F] <= 32'h00058313;
  mem['h0120] <= 32'hf5dff06f;
  mem['h0121] <= 32'h0087e793;
  mem['h0122] <= 32'h00058313;
  mem['h0123] <= 32'hf51ff06f;
  mem['h0124] <= 32'h00058a93;
  mem['h0125] <= 32'h02500793;
  mem['h0126] <= 32'h58f60463;
  mem['h0127] <= 32'h00f50023;
  mem['h0128] <= 32'h000ac783;
  mem['h0129] <= 32'h00150513;
  mem['h012A] <= 32'h56079e63;
  mem['h012B] <= 32'h00050023;
  mem['h012C] <= 32'h03014603;
  mem['h012D] <= 32'hee061ce3;
  mem['h012E] <= 32'h00000513;
  mem['h012F] <= 32'h0400006f;
  mem['h0130] <= 32'h00060893;
  mem['h0131] <= 32'h0015c603;
  mem['h0132] <= 32'h00158a93;
  mem['h0133] <= 32'hfbf60813;
  mem['h0134] <= 32'h0ff87813;
  mem['h0135] <= 32'hfd0c60e3;
  mem['h0136] <= 32'h00001317;
  mem['h0137] <= 32'h8d030313;
  mem['h0138] <= 32'h00281813;
  mem['h0139] <= 32'h00680833;
  mem['h013A] <= 32'h00082803;
  mem['h013B] <= 32'h00680833;
  mem['h013C] <= 32'h00080067;
  mem['h013D] <= 32'h413686b3;
  mem['h013E] <= 32'h00168513;
  mem['h013F] <= 32'h46c12083;
  mem['h0140] <= 32'h46812403;
  mem['h0141] <= 32'h46412483;
  mem['h0142] <= 32'h46012903;
  mem['h0143] <= 32'h45c12983;
  mem['h0144] <= 32'h45812a03;
  mem['h0145] <= 32'h45412a83;
  mem['h0146] <= 32'h45012b03;
  mem['h0147] <= 32'h44c12b83;
  mem['h0148] <= 32'h44812c03;
  mem['h0149] <= 32'h44412c83;
  mem['h014A] <= 32'h44012d03;
  mem['h014B] <= 32'h43c12d83;
  mem['h014C] <= 32'h49010113;
  mem['h014D] <= 32'h00008067;
  mem['h014E] <= 32'h0015c603;
  mem['h014F] <= 32'h00900893;
  mem['h0150] <= 32'h00158813;
  mem['h0151] <= 32'hfd060713;
  mem['h0152] <= 32'h0ff77713;
  mem['h0153] <= 32'h36e8fa63;
  mem['h0154] <= 32'h02a00713;
  mem['h0155] <= 32'h3ae60463;
  mem['h0156] <= 32'h00080593;
  mem['h0157] <= 32'h00000713;
  mem['h0158] <= 32'hec5ff06f;
  mem['h0159] <= 32'h00000693;
  mem['h015A] <= 32'h00900813;
  mem['h015B] <= 32'h00269713;
  mem['h015C] <= 32'h00d70733;
  mem['h015D] <= 32'h00158593;
  mem['h015E] <= 32'h00171713;
  mem['h015F] <= 32'h00c70733;
  mem['h0160] <= 32'h0005c603;
  mem['h0161] <= 32'hfd070693;
  mem['h0162] <= 32'hfd060713;
  mem['h0163] <= 32'h0ff77713;
  mem['h0164] <= 32'hfce87ee3;
  mem['h0165] <= 32'he89ff06f;
  mem['h0166] <= 32'h000a2683;
  mem['h0167] <= 32'h00234603;
  mem['h0168] <= 32'h00230593;
  mem['h0169] <= 32'h004a0a13;
  mem['h016A] <= 32'he606dae3;
  mem['h016B] <= 32'h40d006b3;
  mem['h016C] <= 32'h0107e793;
  mem['h016D] <= 32'he69ff06f;
  mem['h016E] <= 32'h0407e793;
  mem['h016F] <= 32'h06c00713;
  mem['h0170] <= 32'h36e88063;
  mem['h0171] <= 32'h000a2e03;
  mem['h0172] <= 32'h00000593;
  mem['h0173] <= 32'h00000713;
  mem['h0174] <= 32'h00be0633;
  mem['h0175] <= 32'h00064603;
  mem['h0176] <= 32'h00f12423;
  mem['h0177] <= 32'h00d12623;
  mem['h0178] <= 32'h004a0f93;
  mem['h0179] <= 32'h06300393;
  mem['h017A] <= 32'h00000e97;
  mem['h017B] <= 32'h644e8e93;
  mem['h017C] <= 32'h06400b13;
  mem['h017D] <= 32'h00a00b93;
  mem['h017E] <= 32'h03000293;
  mem['h017F] <= 32'h00400313;
  mem['h0180] <= 32'h02e00f13;
  mem['h0181] <= 32'h00170813;
  mem['h0182] <= 32'h04061063;
  mem['h0183] <= 32'h42070793;
  mem['h0184] <= 32'h01010713;
  mem['h0185] <= 32'h00e78733;
  mem['h0186] <= 32'hbe570423;
  mem['h0187] <= 32'h00158593;
  mem['h0188] <= 32'h0a658263;
  mem['h0189] <= 32'h42080793;
  mem['h018A] <= 32'h01010713;
  mem['h018B] <= 32'h00e78633;
  mem['h018C] <= 32'hbfe60423;
  mem['h018D] <= 32'h00be0633;
  mem['h018E] <= 32'h00064603;
  mem['h018F] <= 32'h00180713;
  mem['h0190] <= 32'h00170813;
  mem['h0191] <= 32'hfc0604e3;
  mem['h0192] <= 32'h22c3da63;
  mem['h0193] <= 32'h036667b3;
  mem['h0194] <= 32'h42070693;
  mem['h0195] <= 32'h01010893;
  mem['h0196] <= 32'h011688b3;
  mem['h0197] <= 32'h00088693;
  mem['h0198] <= 32'h42080813;
  mem['h0199] <= 32'h01010893;
  mem['h019A] <= 32'h01180833;
  mem['h019B] <= 32'h01012223;
  mem['h019C] <= 32'h00270713;
  mem['h019D] <= 32'h000e8893;
  mem['h019E] <= 32'h00170813;
  mem['h019F] <= 32'h03664633;
  mem['h01A0] <= 32'h0377ca33;
  mem['h01A1] <= 32'h00ce8633;
  mem['h01A2] <= 32'h00064603;
  mem['h01A3] <= 32'hbec68423;
  mem['h01A4] <= 32'h014e8a33;
  mem['h01A5] <= 32'h0377e633;
  mem['h01A6] <= 32'h000a4a03;
  mem['h01A7] <= 32'h00412783;
  mem['h01A8] <= 32'hbf478423;
  mem['h01A9] <= 32'h00c888b3;
  mem['h01AA] <= 32'h0008c603;
  mem['h01AB] <= 32'h42070793;
  mem['h01AC] <= 32'h01010713;
  mem['h01AD] <= 32'h00e78733;
  mem['h01AE] <= 32'hbec70423;
  mem['h01AF] <= 32'h00158593;
  mem['h01B0] <= 32'hf66592e3;
  mem['h01B1] <= 32'h00812783;
  mem['h01B2] <= 32'h00c12683;
  mem['h01B3] <= 32'h0107f793;
  mem['h01B4] <= 32'h02079663;
  mem['h01B5] <= 32'hfff68613;
  mem['h01B6] <= 32'h4ad85e63;
  mem['h01B7] <= 32'h410687b3;
  mem['h01B8] <= 32'h00f507b3;
  mem['h01B9] <= 32'h02000713;
  mem['h01BA] <= 32'h00150513;
  mem['h01BB] <= 32'hfee50fa3;
  mem['h01BC] <= 32'hfea79ce3;
  mem['h01BD] <= 32'h40d806b3;
  mem['h01BE] <= 32'h00c686b3;
  mem['h01BF] <= 32'h01810613;
  mem['h01C0] <= 32'h010507b3;
  mem['h01C1] <= 32'h00050713;
  mem['h01C2] <= 32'h00064583;
  mem['h01C3] <= 32'h00170713;
  mem['h01C4] <= 32'h00160613;
  mem['h01C5] <= 32'hfeb70fa3;
  mem['h01C6] <= 32'hfee798e3;
  mem['h01C7] <= 32'h44d85863;
  mem['h01C8] <= 32'h00d50533;
  mem['h01C9] <= 32'h02000713;
  mem['h01CA] <= 32'h00178793;
  mem['h01CB] <= 32'hfee78fa3;
  mem['h01CC] <= 32'hfea79ce3;
  mem['h01CD] <= 32'h001ac783;
  mem['h01CE] <= 32'h001a8313;
  mem['h01CF] <= 32'h000f8a13;
  mem['h01D0] <= 32'hc40794e3;
  mem['h01D1] <= 32'hc5dff06f;
  mem['h01D2] <= 32'h0407e793;
  mem['h01D3] <= 32'h01000613;
  mem['h01D4] <= 32'h004a0813;
  mem['h01D5] <= 32'h000a2583;
  mem['h01D6] <= 32'h00080a13;
  mem['h01D7] <= 32'h909ff0ef;
  mem['h01D8] <= 32'h001ac783;
  mem['h01D9] <= 32'h001a8313;
  mem['h01DA] <= 32'hc20790e3;
  mem['h01DB] <= 32'hc35ff06f;
  mem['h01DC] <= 32'h00058a93;
  mem['h01DD] <= 32'h0107f793;
  mem['h01DE] <= 32'h004a0613;
  mem['h01DF] <= 32'h001a8313;
  mem['h01E0] <= 32'h2c078a63;
  mem['h01E1] <= 32'h000a2783;
  mem['h01E2] <= 32'h00100593;
  mem['h01E3] <= 32'h00150713;
  mem['h01E4] <= 32'h00f50023;
  mem['h01E5] <= 32'h02000793;
  mem['h01E6] <= 32'h00d50533;
  mem['h01E7] <= 32'h40d5d463;
  mem['h01E8] <= 32'h00170713;
  mem['h01E9] <= 32'hfef70fa3;
  mem['h01EA] <= 32'hfea71ce3;
  mem['h01EB] <= 32'h001ac783;
  mem['h01EC] <= 32'h00060a13;
  mem['h01ED] <= 32'hbc079ae3;
  mem['h01EE] <= 32'hbe9ff06f;
  mem['h01EF] <= 32'h00058a93;
  mem['h01F0] <= 32'h000a2603;
  mem['h01F1] <= 32'h004a0a13;
  mem['h01F2] <= 32'h28060063;
  mem['h01F3] <= 32'h00064583;
  mem['h01F4] <= 32'h30058e63;
  mem['h01F5] <= 32'h30070c63;
  mem['h01F6] <= 32'h00060593;
  mem['h01F7] <= 32'h00c0006f;
  mem['h01F8] <= 32'h40e58833;
  mem['h01F9] <= 32'h00c80863;
  mem['h01FA] <= 32'h0015c803;
  mem['h01FB] <= 32'h00158593;
  mem['h01FC] <= 32'hfe0818e3;
  mem['h01FD] <= 32'h0107f713;
  mem['h01FE] <= 32'h40c587b3;
  mem['h01FF] <= 32'h28070c63;
  mem['h0200] <= 32'h3af05c63;
  mem['h0201] <= 32'h00f60833;
  mem['h0202] <= 32'h00050713;
  mem['h0203] <= 32'h00064583;
  mem['h0204] <= 32'h00160613;
  mem['h0205] <= 32'h00170713;
  mem['h0206] <= 32'hfeb70fa3;
  mem['h0207] <= 32'hff0618e3;
  mem['h0208] <= 32'h00f50733;
  mem['h0209] <= 32'h40f68533;
  mem['h020A] <= 32'h001a8313;
  mem['h020B] <= 32'h00a70533;
  mem['h020C] <= 32'h02000613;
  mem['h020D] <= 32'h34d7d863;
  mem['h020E] <= 32'h00170713;
  mem['h020F] <= 32'hfec70fa3;
  mem['h0210] <= 32'hfea71ce3;
  mem['h0211] <= 32'h001ac783;
  mem['h0212] <= 32'hb40790e3;
  mem['h0213] <= 32'hb55ff06f;
  mem['h0214] <= 32'h00058a93;
  mem['h0215] <= 32'hfff00613;
  mem['h0216] <= 32'h1ec68263;
  mem['h0217] <= 32'h000a2583;
  mem['h0218] <= 32'h01000613;
  mem['h0219] <= 32'h004a0a13;
  mem['h021A] <= 32'hffcff0ef;
  mem['h021B] <= 32'h001ac783;
  mem['h021C] <= 32'h001a8313;
  mem['h021D] <= 32'hb0079ae3;
  mem['h021E] <= 32'hb29ff06f;
  mem['h021F] <= 32'h00900793;
  mem['h0220] <= 32'h000e8893;
  mem['h0221] <= 32'he2c7d0e3;
  mem['h0222] <= 32'h00a00a13;
  mem['h0223] <= 32'h034647b3;
  mem['h0224] <= 32'h00000897;
  mem['h0225] <= 32'h39c88893;
  mem['h0226] <= 32'h42070713;
  mem['h0227] <= 32'h01010693;
  mem['h0228] <= 32'h00d706b3;
  mem['h0229] <= 32'h00080713;
  mem['h022A] <= 32'h00180813;
  mem['h022B] <= 32'h03466633;
  mem['h022C] <= 32'h00f88a33;
  mem['h022D] <= 32'h000a4a03;
  mem['h022E] <= 32'hbf468423;
  mem['h022F] <= 32'hde9ff06f;
  mem['h0230] <= 32'h00000713;
  mem['h0231] <= 32'h00070313;
  mem['h0232] <= 32'h00231713;
  mem['h0233] <= 32'h00670733;
  mem['h0234] <= 32'h00180813;
  mem['h0235] <= 32'h00171713;
  mem['h0236] <= 32'h00c70733;
  mem['h0237] <= 32'h00084603;
  mem['h0238] <= 32'hfd070313;
  mem['h0239] <= 32'hfd060593;
  mem['h023A] <= 32'h0ff5f593;
  mem['h023B] <= 32'hfcb8fee3;
  mem['h023C] <= 32'h00030713;
  mem['h023D] <= 32'h00080593;
  mem['h023E] <= 32'hb2dff06f;
  mem['h023F] <= 32'h000a2703;
  mem['h0240] <= 32'h00258813;
  mem['h0241] <= 32'h0025c603;
  mem['h0242] <= 32'hfff74593;
  mem['h0243] <= 32'h41f5d593;
  mem['h0244] <= 32'h00b77733;
  mem['h0245] <= 32'h004a0a13;
  mem['h0246] <= 32'h00080593;
  mem['h0247] <= 32'hb09ff06f;
  mem['h0248] <= 32'h0407f713;
  mem['h0249] <= 32'h00000317;
  mem['h024A] <= 32'h30830313;
  mem['h024B] <= 32'h00070663;
  mem['h024C] <= 32'h00000317;
  mem['h024D] <= 32'h32430313;
  mem['h024E] <= 32'h000a2e83;
  mem['h024F] <= 32'h00000613;
  mem['h0250] <= 32'h00000893;
  mem['h0251] <= 32'h00600e13;
  mem['h0252] <= 32'h03a00f13;
  mem['h0253] <= 32'h0140006f;
  mem['h0254] <= 32'h42288713;
  mem['h0255] <= 32'h00770833;
  mem['h0256] <= 32'h00388893;
  mem['h0257] <= 32'hbfe80423;
  mem['h0258] <= 32'h00ce8733;
  mem['h0259] <= 32'h00074703;
  mem['h025A] <= 32'h01010393;
  mem['h025B] <= 32'h00160613;
  mem['h025C] <= 32'h00475813;
  mem['h025D] <= 32'h00f77713;
  mem['h025E] <= 32'h00e30733;
  mem['h025F] <= 32'h01030833;
  mem['h0260] <= 32'h00074f83;
  mem['h0261] <= 32'h00084283;
  mem['h0262] <= 32'h42088713;
  mem['h0263] <= 32'h00770733;
  mem['h0264] <= 32'hbe570423;
  mem['h0265] <= 32'hbff704a3;
  mem['h0266] <= 32'hfbc61ce3;
  mem['h0267] <= 32'h0107f793;
  mem['h0268] <= 32'h02079863;
  mem['h0269] <= 32'h01100793;
  mem['h026A] <= 32'hfff68613;
  mem['h026B] <= 32'h20d7de63;
  mem['h026C] <= 32'hfef68793;
  mem['h026D] <= 32'h00f507b3;
  mem['h026E] <= 32'h02000713;
  mem['h026F] <= 32'h00150513;
  mem['h0270] <= 32'hfee50fa3;
  mem['h0271] <= 32'hfea79ce3;
  mem['h0272] <= 32'h40d60633;
  mem['h0273] <= 32'h01160693;
  mem['h0274] <= 32'h01810613;
  mem['h0275] <= 32'h01150793;
  mem['h0276] <= 32'h00050713;
  mem['h0277] <= 32'h00064803;
  mem['h0278] <= 32'h00170713;
  mem['h0279] <= 32'h00160613;
  mem['h027A] <= 32'hff070fa3;
  mem['h027B] <= 32'hfef718e3;
  mem['h027C] <= 32'h01100613;
  mem['h027D] <= 32'h1ad65463;
  mem['h027E] <= 32'h00d50533;
  mem['h027F] <= 32'h02000713;
  mem['h0280] <= 32'h00178793;
  mem['h0281] <= 32'hfee78fa3;
  mem['h0282] <= 32'hfef51ce3;
  mem['h0283] <= 32'h0025c783;
  mem['h0284] <= 32'h004a0a13;
  mem['h0285] <= 32'h00258313;
  mem['h0286] <= 32'h960798e3;
  mem['h0287] <= 32'h985ff06f;
  mem['h0288] <= 32'h000ac783;
  mem['h0289] <= 32'h00f50023;
  mem['h028A] <= 32'h001ac783;
  mem['h028B] <= 32'h00150513;
  mem['h028C] <= 32'h001a8313;
  mem['h028D] <= 32'h94079ae3;
  mem['h028E] <= 32'h969ff06f;
  mem['h028F] <= 32'h0017e793;
  mem['h0290] <= 32'h00800693;
  mem['h0291] <= 32'he19ff06f;
  mem['h0292] <= 32'h00000617;
  mem['h0293] <= 32'h23460613;
  mem['h0294] <= 32'hd85ff06f;
  mem['h0295] <= 32'h00100793;
  mem['h0296] <= 32'h0ed7dc63;
  mem['h0297] <= 32'hfff68793;
  mem['h0298] <= 32'h00f507b3;
  mem['h0299] <= 32'h02000713;
  mem['h029A] <= 32'h00150513;
  mem['h029B] <= 32'hfee50fa3;
  mem['h029C] <= 32'hfef51ce3;
  mem['h029D] <= 32'h00000693;
  mem['h029E] <= 32'hd0dff06f;
  mem['h029F] <= 32'h0027e793;
  mem['h02A0] <= 32'h00a00613;
  mem['h02A1] <= 32'hccdff06f;
  mem['h02A2] <= 32'h03010993;
  mem['h02A3] <= 32'h00098513;
  mem['h02A4] <= 32'h911ff06f;
  mem['h02A5] <= 32'hfff68813;
  mem['h02A6] <= 32'h12d7d463;
  mem['h02A7] <= 32'h40f68733;
  mem['h02A8] <= 32'h00e50733;
  mem['h02A9] <= 32'h02000593;
  mem['h02AA] <= 32'h00150513;
  mem['h02AB] <= 32'hfeb50fa3;
  mem['h02AC] <= 32'hfee51ce3;
  mem['h02AD] <= 32'h40d786b3;
  mem['h02AE] <= 32'h010686b3;
  mem['h02AF] <= 32'hd45ff06f;
  mem['h02B0] <= 32'h0027e793;
  mem['h02B1] <= 32'h004a0813;
  mem['h02B2] <= 32'h00058a93;
  mem['h02B3] <= 32'h00a00613;
  mem['h02B4] <= 32'hc85ff06f;
  mem['h02B5] <= 32'h00800613;
  mem['h02B6] <= 32'hc79ff06f;
  mem['h02B7] <= 32'h00a00613;
  mem['h02B8] <= 32'hc71ff06f;
  mem['h02B9] <= 32'h00058a93;
  mem['h02BA] <= 32'haddff06f;
  mem['h02BB] <= 32'h0107f793;
  mem['h02BC] <= 32'h08078263;
  mem['h02BD] <= 32'h00050713;
  mem['h02BE] <= 32'h00000793;
  mem['h02BF] <= 32'hd29ff06f;
  mem['h02C0] <= 32'h0407e793;
  mem['h02C1] <= 32'h00058a93;
  mem['h02C2] <= 32'habdff06f;
  mem['h02C3] <= 32'h004a0813;
  mem['h02C4] <= 32'h00058a93;
  mem['h02C5] <= 32'h00a00613;
  mem['h02C6] <= 32'hc3dff06f;
  mem['h02C7] <= 32'h0407e793;
  mem['h02C8] <= 32'h004a0813;
  mem['h02C9] <= 32'h00058a93;
  mem['h02CA] <= 32'h01000613;
  mem['h02CB] <= 32'hc29ff06f;
  mem['h02CC] <= 32'h004a0813;
  mem['h02CD] <= 32'h00058a93;
  mem['h02CE] <= 32'h01000613;
  mem['h02CF] <= 32'hc19ff06f;
  mem['h02D0] <= 32'h004a0813;
  mem['h02D1] <= 32'h00058a93;
  mem['h02D2] <= 32'h00800613;
  mem['h02D3] <= 32'hc09ff06f;
  mem['h02D4] <= 32'h000a2783;
  mem['h02D5] <= 32'h00150513;
  mem['h02D6] <= 32'h00060a13;
  mem['h02D7] <= 32'hfef50fa3;
  mem['h02D8] <= 32'h001ac783;
  mem['h02D9] <= 32'h820792e3;
  mem['h02DA] <= 32'h839ff06f;
  mem['h02DB] <= 32'h00078513;
  mem['h02DC] <= 32'hbc5ff06f;
  mem['h02DD] <= 32'hfff68813;
  mem['h02DE] <= 32'hf2d042e3;
  mem['h02DF] <= 32'h001a8313;
  mem['h02E0] <= 32'h00050713;
  mem['h02E1] <= 32'h001ac783;
  mem['h02E2] <= 32'h00070513;
  mem['h02E3] <= 32'hfe079e63;
  mem['h02E4] <= 32'h811ff06f;
  mem['h02E5] <= 32'h00060693;
  mem['h02E6] <= 32'hb65ff06f;
  mem['h02E7] <= 32'h00070513;
  mem['h02E8] <= 32'he6dff06f;
  mem['h02E9] <= 32'h001ac783;
  mem['h02EA] <= 32'h00060a13;
  mem['h02EB] <= 32'h00070513;
  mem['h02EC] <= 32'hfc079c63;
  mem['h02ED] <= 32'hfecff06f;
  mem['h02EE] <= 32'h00050713;
  mem['h02EF] <= 32'hc69ff06f;
  mem['h02F0] <= 32'h00080693;
  mem['h02F1] <= 32'hc3dff06f;
  mem['h02F2] <= 32'h00060693;
  mem['h02F3] <= 32'he05ff06f;
  mem['h02F4] <= 32'h200007b7;
  mem['h02F5] <= 32'h0007a703;
  mem['h02F6] <= 32'h00176713;
  mem['h02F7] <= 32'h00e7a023;
  mem['h02F8] <= 32'h0007a703;
  mem['h02F9] <= 32'h00276713;
  mem['h02FA] <= 32'h00e7a023;
  mem['h02FB] <= 32'h43d00713;
  mem['h02FC] <= 32'h00e79123;
  mem['h02FD] <= 32'h00008067;
  mem['h02FE] <= 32'h20000737;
  mem['h02FF] <= 32'h00472783;
  mem['h0300] <= 32'h0037d793;
  mem['h0301] <= 32'h0017f793;
  mem['h0302] <= 32'hfe079ae3;
  mem['h0303] <= 32'h00874503;
  mem['h0304] <= 32'h00008067;
  mem['h0305] <= 32'h6c6c6568;
  mem['h0306] <= 32'h0000006f;
  mem['h0307] <= 32'h656e6f64;
  mem['h0308] <= 32'h00000000;
  mem['h0309] <= 32'h00000066;
  mem['h030A] <= 32'h00006325;
  mem['h030B] <= 32'h33323130;
  mem['h030C] <= 32'h37363534;
  mem['h030D] <= 32'h62613938;
  mem['h030E] <= 32'h66656463;
  mem['h030F] <= 32'h6a696867;
  mem['h0310] <= 32'h6e6d6c6b;
  mem['h0311] <= 32'h7271706f;
  mem['h0312] <= 32'h76757473;
  mem['h0313] <= 32'h7a797877;
  mem['h0314] <= 32'h00000000;
  mem['h0315] <= 32'h33323130;
  mem['h0316] <= 32'h37363534;
  mem['h0317] <= 32'h42413938;
  mem['h0318] <= 32'h46454443;
  mem['h0319] <= 32'h4a494847;
  mem['h031A] <= 32'h4e4d4c4b;
  mem['h031B] <= 32'h5251504f;
  mem['h031C] <= 32'h56555453;
  mem['h031D] <= 32'h5a595857;
  mem['h031E] <= 32'h00000000;
  mem['h031F] <= 32'h4c554e3c;
  mem['h0320] <= 32'h00003e4c;
  mem['h0321] <= 32'hfffff800;
  mem['h0322] <= 32'hfffff780;
  mem['h0323] <= 32'hfffff780;
  mem['h0324] <= 32'hfffff7f4;
  mem['h0325] <= 32'hfffff780;
  mem['h0326] <= 32'hfffff780;
  mem['h0327] <= 32'hfffff780;
  mem['h0328] <= 32'hfffff780;
  mem['h0329] <= 32'hfffff780;
  mem['h032A] <= 32'hfffff780;
  mem['h032B] <= 32'hfffff780;
  mem['h032C] <= 32'hfffff7e8;
  mem['h032D] <= 32'hfffff780;
  mem['h032E] <= 32'hfffff7dc;
  mem['h032F] <= 32'hfffff780;
  mem['h0330] <= 32'hfffff780;
  mem['h0331] <= 32'hfffff7d0;
  mem['h0332] <= 32'hfffffe38;
  mem['h0333] <= 32'hfffff7c8;
  mem['h0334] <= 32'hfffff7c8;
  mem['h0335] <= 32'hfffff7c8;
  mem['h0336] <= 32'hfffff7c8;
  mem['h0337] <= 32'hfffff7c8;
  mem['h0338] <= 32'hfffff7c8;
  mem['h0339] <= 32'hfffff7c8;
  mem['h033A] <= 32'hfffff7c8;
  mem['h033B] <= 32'hfffff7c8;
  mem['h033C] <= 32'hfffff7c8;
  mem['h033D] <= 32'hfffff7c8;
  mem['h033E] <= 32'hfffff7c8;
  mem['h033F] <= 32'hfffff7c8;
  mem['h0340] <= 32'hfffff7c8;
  mem['h0341] <= 32'hfffff7c8;
  mem['h0342] <= 32'hfffff7c8;
  mem['h0343] <= 32'hfffff7c8;
  mem['h0344] <= 32'hfffff7c8;
  mem['h0345] <= 32'hfffff7c8;
  mem['h0346] <= 32'hfffff7c8;
  mem['h0347] <= 32'hfffff7c8;
  mem['h0348] <= 32'hfffff7c8;
  mem['h0349] <= 32'hfffffe54;
  mem['h034A] <= 32'hfffff7c8;
  mem['h034B] <= 32'hfffff7c8;
  mem['h034C] <= 32'hfffff7c8;
  mem['h034D] <= 32'hfffff7c8;
  mem['h034E] <= 32'hfffff7c8;
  mem['h034F] <= 32'hfffff7c8;
  mem['h0350] <= 32'hfffff7c8;
  mem['h0351] <= 32'hfffff7c8;
  mem['h0352] <= 32'hfffffe1c;
  mem['h0353] <= 32'hfffff7c8;
  mem['h0354] <= 32'hfffffaa8;
  mem['h0355] <= 32'hfffffdf8;
  mem['h0356] <= 32'hfffff7c8;
  mem['h0357] <= 32'hfffff7c8;
  mem['h0358] <= 32'hfffff7c8;
  mem['h0359] <= 32'hfffff7c8;
  mem['h035A] <= 32'hfffffdf8;
  mem['h035B] <= 32'hfffff7c8;
  mem['h035C] <= 32'hfffff7c8;
  mem['h035D] <= 32'hfffff7c8;
  mem['h035E] <= 32'hfffff7c8;
  mem['h035F] <= 32'hfffff7c8;
  mem['h0360] <= 32'hfffffe78;
  mem['h0361] <= 32'hfffffb88;
  mem['h0362] <= 32'hfffff7c8;
  mem['h0363] <= 32'hfffff7c8;
  mem['h0364] <= 32'hfffffaf4;
  mem['h0365] <= 32'hfffff7c8;
  mem['h0366] <= 32'hfffffe44;
  mem['h0367] <= 32'hfffff7c8;
  mem['h0368] <= 32'hfffff7c8;
  mem['h0369] <= 32'hfffffe68;
  mem['h036A] <= 32'hfffff810;
  mem['h036B] <= 32'hfffff6ec;
  mem['h036C] <= 32'hfffff6ec;
  mem['h036D] <= 32'hfffff6ec;
  mem['h036E] <= 32'hfffff6ec;
  mem['h036F] <= 32'hfffff6ec;
  mem['h0370] <= 32'hfffff6ec;
  mem['h0371] <= 32'hfffff6ec;
  mem['h0372] <= 32'hfffff6ec;
  mem['h0373] <= 32'hfffff6ec;
  mem['h0374] <= 32'hfffff6ec;
  mem['h0375] <= 32'hfffff6ec;
  mem['h0376] <= 32'hfffff6ec;
  mem['h0377] <= 32'hfffff6ec;
  mem['h0378] <= 32'hfffff6ec;
  mem['h0379] <= 32'hfffff6ec;
  mem['h037A] <= 32'hfffff6ec;
  mem['h037B] <= 32'hfffff6ec;
  mem['h037C] <= 32'hfffff6ec;
  mem['h037D] <= 32'hfffff6ec;
  mem['h037E] <= 32'hfffff6ec;
  mem['h037F] <= 32'hfffff6ec;
  mem['h0380] <= 32'hfffff6ec;
  mem['h0381] <= 32'hfffff9a0;
  mem['h0382] <= 32'hfffff6ec;
  mem['h0383] <= 32'hfffff6ec;
  mem['h0384] <= 32'hfffff6ec;
  mem['h0385] <= 32'hfffff6ec;
  mem['h0386] <= 32'hfffff6ec;
  mem['h0387] <= 32'hfffff6ec;
  mem['h0388] <= 32'hfffff6ec;
  mem['h0389] <= 32'hfffff6ec;
  mem['h038A] <= 32'hfffff814;
  mem['h038B] <= 32'hfffff6ec;
  mem['h038C] <= 32'hfffff9cc;
  mem['h038D] <= 32'hfffffcd4;
  mem['h038E] <= 32'hfffff6ec;
  mem['h038F] <= 32'hfffff6ec;
  mem['h0390] <= 32'hfffff6ec;
  mem['h0391] <= 32'hfffff6ec;
  mem['h0392] <= 32'hfffffcd4;
  mem['h0393] <= 32'hfffff6ec;
  mem['h0394] <= 32'hfffff6ec;
  mem['h0395] <= 32'hfffff6ec;
  mem['h0396] <= 32'hfffff6ec;
  mem['h0397] <= 32'hfffff6ec;
  mem['h0398] <= 32'hfffffd2c;
  mem['h0399] <= 32'hfffffaac;
  mem['h039A] <= 32'hfffff6ec;
  mem['h039B] <= 32'hfffff6ec;
  mem['h039C] <= 32'hfffffa18;
  mem['h039D] <= 32'hfffff6ec;
  mem['h039E] <= 32'hfffffd34;
  mem['h039F] <= 32'hfffff6ec;
  mem['h03A0] <= 32'hfffff6ec;
  mem['h03A1] <= 32'hfffff9a4;

  end

  always @(posedge clk) mem_data <= mem[mem_addr];

  // ============================================================================

  reg o_ready;

  always @(posedge clk or negedge rstn)
    if (!rstn) o_ready <= 1'd0;
    else o_ready <= valid && ((addr & MEM_ADDR_MASK) != 0);

  // Output connectins
  assign ready    = o_ready;
  assign rdata    = mem_data;
  assign mem_addr = addr[MEM_SIZE_BITS+1:2];

endmodule

