// coz_yazmacoku.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module coz_yazmacoku(
    input clk_i,
    input rst_i


);


endmodule
