
module RAM256x8 (CLK,
    EN0,
    WE0,
    A0,
    Di0,
    Do0);
 input CLK;
 input EN0;
 input WE0;
 input [7:0] A0;
 input [7:0] Di0;
 output [7:0] Do0;

 wire \BANK128[0].RAM128.A0BUF[0].X ;
 wire \BANK128[0].RAM128.A0BUF[1].X ;
 wire \BANK128[0].RAM128.A0BUF[2].X ;
 wire \BANK128[0].RAM128.A0BUF[3].X ;
 wire \BANK128[0].RAM128.A0BUF[4].X ;
 wire \BANK128[0].RAM128.A0BUF[5].X ;
 wire \BANK128[0].RAM128.A0BUF[6].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[4].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].A ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].A ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].A ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].A ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].A ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].A ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].A ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].A ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.Do0[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.EN0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.EN0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.WE0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.EN0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[0].RAM32.WE0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[4].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.Do0[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.EN0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.EN0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.WE0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.EN0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[4].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.Do0[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.EN0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.EN0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.WE0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.EN0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[4].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.Do0[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.EN0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.EN0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.WE0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.EN0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[0].RAM128.DEC0.EN ;
 wire \BANK128[0].RAM128.Do0MUX.SEL0 ;
 wire \BANK128[0].RAM128.Do0MUX.SEL1 ;
 wire \BANK128[0].RAM128.Do0[0] ;
 wire \BANK128[0].RAM128.Do0[1] ;
 wire \BANK128[0].RAM128.Do0[2] ;
 wire \BANK128[0].RAM128.Do0[3] ;
 wire \BANK128[0].RAM128.Do0[4] ;
 wire \BANK128[0].RAM128.Do0[5] ;
 wire \BANK128[0].RAM128.Do0[6] ;
 wire \BANK128[0].RAM128.Do0[7] ;
 wire \BANK128[0].RAM128.EN0 ;
 wire \BANK128[1].RAM128.A0BUF[0].X ;
 wire \BANK128[1].RAM128.A0BUF[1].X ;
 wire \BANK128[1].RAM128.A0BUF[2].X ;
 wire \BANK128[1].RAM128.A0BUF[3].X ;
 wire \BANK128[1].RAM128.A0BUF[4].X ;
 wire \BANK128[1].RAM128.A0BUF[5].X ;
 wire \BANK128[1].RAM128.A0BUF[6].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[4].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].A ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].A ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].A ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].A ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].A ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].A ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].A ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].A ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.Do0[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.EN0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.EN0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.WE0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.EN0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[0].RAM32.WE0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[4].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.Do0[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.EN0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.EN0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.WE0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.EN0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[4].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.Do0[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.EN0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.EN0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.WE0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.EN0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[4].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.Do0[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.EN0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.EN0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.WE0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.EN0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BANK128[1].RAM128.DEC0.EN ;
 wire \BANK128[1].RAM128.Do0MUX.SEL0 ;
 wire \BANK128[1].RAM128.Do0MUX.SEL1 ;
 wire \BANK128[1].RAM128.Do0[0] ;
 wire \BANK128[1].RAM128.Do0[1] ;
 wire \BANK128[1].RAM128.Do0[2] ;
 wire \BANK128[1].RAM128.Do0[3] ;
 wire \BANK128[1].RAM128.Do0[4] ;
 wire \BANK128[1].RAM128.Do0[5] ;
 wire \BANK128[1].RAM128.Do0[6] ;
 wire \BANK128[1].RAM128.Do0[7] ;
 wire \BANK128[1].RAM128.EN0 ;
 wire \Do0MUX.SEL ;

 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.A0BUF[0].__cell__  (.A(A0[0]),
    .X(\BANK128[0].RAM128.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.A0BUF[1].__cell__  (.A(A0[1]),
    .X(\BANK128[0].RAM128.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.A0BUF[2].__cell__  (.A(A0[2]),
    .X(\BANK128[0].RAM128.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.A0BUF[3].__cell__  (.A(A0[3]),
    .X(\BANK128[0].RAM128.A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.A0BUF[4].__cell__  (.A(A0[4]),
    .X(\BANK128[0].RAM128.A0BUF[4].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.A0BUF[5].__cell__  (.A(A0[5]),
    .X(\BANK128[0].RAM128.A0BUF[5].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.A0BUF[6].__cell__  (.A(A0[6]),
    .X(\BANK128[0].RAM128.A0BUF[6].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[0].__cell__  (.A(\BANK128[0].RAM128.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[1].__cell__  (.A(\BANK128[0].RAM128.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[2].__cell__  (.A(\BANK128[0].RAM128.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[3].__cell__  (.A(\BANK128[0].RAM128.A0BUF[3].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[4].__cell__  (.A(\BANK128[0].RAM128.A0BUF[4].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[4].X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.DEC0.AND0  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[4].X ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.EN0 ));
 sky130_fd_sc_hd__and2_2 \BANK128[0].RAM128.BLOCK[0].RAM32.DEC0.AND1  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[4].X ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.EN0 ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].A ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].A ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].A ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].A ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].A ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].A ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].A ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].A ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[0]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[0] ),
    .A1(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[0] ),
    .S(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[0] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[1]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[1] ),
    .A1(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[1] ),
    .S(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[1] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[2]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[2] ),
    .A1(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[2] ),
    .S(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[2] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[3]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[3] ),
    .A1(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[3] ),
    .S(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[3] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[4]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[4] ),
    .A1(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[4] ),
    .S(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[4] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[5]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[5] ),
    .A1(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[5] ),
    .S(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[5] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[6]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[6] ),
    .A1(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[6] ),
    .S(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[6] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[7]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[7] ),
    .A1(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[7] ),
    .S(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[7] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.SEL0BUF[0]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[4].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.EN0BUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[3].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.DEC0.AND0  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.DEC0.AND1  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.EN0BUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.TIE0[0].__cell__  (.LO(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.A0BUF[3].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.DEC0.AND0  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.DEC0.AND1  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.EN0BUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.TIE0[0].__cell__  (.LO(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[0].RAM32.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[0].__cell__  (.A(\BANK128[0].RAM128.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[1].__cell__  (.A(\BANK128[0].RAM128.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[2].__cell__  (.A(\BANK128[0].RAM128.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[3].__cell__  (.A(\BANK128[0].RAM128.A0BUF[3].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[4].__cell__  (.A(\BANK128[0].RAM128.A0BUF[4].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[4].X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.DEC0.AND0  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[4].X ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.EN0 ));
 sky130_fd_sc_hd__and2_2 \BANK128[0].RAM128.BLOCK[1].RAM32.DEC0.AND1  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[4].X ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.EN0 ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].A ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].A ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].A ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].A ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].A ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].A ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].A ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].A ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[0]  (.A0(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[0] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[0] ),
    .S(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[0] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[1]  (.A0(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[1] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[1] ),
    .S(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[1] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[2]  (.A0(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[2] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[2] ),
    .S(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[2] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[3]  (.A0(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[3] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[3] ),
    .S(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[3] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[4]  (.A0(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[4] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[4] ),
    .S(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[4] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[5]  (.A0(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[5] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[5] ),
    .S(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[5] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[6]  (.A0(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[6] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[6] ),
    .S(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[6] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[7]  (.A0(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[7] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[7] ),
    .S(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[7] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.SEL0BUF[0]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[4].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.EN0BUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[3].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.DEC0.AND0  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.DEC0.AND1  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.EN0BUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.TIE0[0].__cell__  (.LO(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.A0BUF[3].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.DEC0.AND0  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.DEC0.AND1  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.EN0BUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.TIE0[0].__cell__  (.LO(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[1].RAM32.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[0].__cell__  (.A(\BANK128[0].RAM128.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[1].__cell__  (.A(\BANK128[0].RAM128.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[2].__cell__  (.A(\BANK128[0].RAM128.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[3].__cell__  (.A(\BANK128[0].RAM128.A0BUF[3].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[4].__cell__  (.A(\BANK128[0].RAM128.A0BUF[4].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[4].X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.DEC0.AND0  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[4].X ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.EN0 ));
 sky130_fd_sc_hd__and2_2 \BANK128[0].RAM128.BLOCK[2].RAM32.DEC0.AND1  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[4].X ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.EN0 ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].A ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].A ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].A ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].A ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].A ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].A ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].A ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].A ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[0]  (.A0(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[0] ),
    .A1(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[0] ),
    .S(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[0] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[1]  (.A0(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[1] ),
    .A1(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[1] ),
    .S(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[1] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[2]  (.A0(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[2] ),
    .A1(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[2] ),
    .S(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[2] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[3]  (.A0(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[3] ),
    .A1(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[3] ),
    .S(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[3] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[4]  (.A0(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[4] ),
    .A1(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[4] ),
    .S(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[4] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[5]  (.A0(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[5] ),
    .A1(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[5] ),
    .S(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[5] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[6]  (.A0(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[6] ),
    .A1(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[6] ),
    .S(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[6] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[7]  (.A0(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[7] ),
    .A1(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[7] ),
    .S(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[7] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.SEL0BUF[0]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[4].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.EN0BUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[3].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.DEC0.AND0  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.DEC0.AND1  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.EN0BUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.TIE0[0].__cell__  (.LO(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.A0BUF[3].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.DEC0.AND0  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.DEC0.AND1  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.EN0BUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.TIE0[0].__cell__  (.LO(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[2].RAM32.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[0].__cell__  (.A(\BANK128[0].RAM128.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[1].__cell__  (.A(\BANK128[0].RAM128.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[2].__cell__  (.A(\BANK128[0].RAM128.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[3].__cell__  (.A(\BANK128[0].RAM128.A0BUF[3].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[4].__cell__  (.A(\BANK128[0].RAM128.A0BUF[4].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[4].X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.DEC0.AND0  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[4].X ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.EN0 ));
 sky130_fd_sc_hd__and2_2 \BANK128[0].RAM128.BLOCK[3].RAM32.DEC0.AND1  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[4].X ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.EN0 ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].A ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].A ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].A ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].A ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].A ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].A ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].A ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].A ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[0]  (.A0(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[0] ),
    .A1(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[0] ),
    .S(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[0] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[1]  (.A0(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[1] ),
    .A1(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[1] ),
    .S(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[1] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[2]  (.A0(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[2] ),
    .A1(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[2] ),
    .S(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[2] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[3]  (.A0(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[3] ),
    .A1(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[3] ),
    .S(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[3] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[4]  (.A0(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[4] ),
    .A1(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[4] ),
    .S(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[4] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[5]  (.A0(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[5] ),
    .A1(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[5] ),
    .S(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[5] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[6]  (.A0(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[6] ),
    .A1(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[6] ),
    .S(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[6] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[7]  (.A0(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[7] ),
    .A1(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[7] ),
    .S(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[7] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.SEL0BUF[0]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[4].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.EN0BUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[3].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.DEC0.AND0  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.DEC0.AND1  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.EN0BUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.TIE0[0].__cell__  (.LO(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.A0BUF[3].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.DEC0.AND0  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.DEC0.AND1  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.EN0BUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[0].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.TIE0[0].__cell__  (.LO(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.BLOCK[3].RAM32.WEBUF[0].__cell__  (.A(\BANK128[0].RAM128.BLOCK[0].RAM32.WE0 ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.WE0 ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[0].RAM128.CLKBUF.__cell__  (.A(CLK),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.CLK ));
 sky130_fd_sc_hd__nor3b_2 \BANK128[0].RAM128.DEC0.AND0  (.A(\BANK128[0].RAM128.A0BUF[5].X ),
    .B(\BANK128[0].RAM128.A0BUF[6].X ),
    .C_N(\BANK128[0].RAM128.DEC0.EN ),
    .Y(\BANK128[0].RAM128.BLOCK[0].RAM32.EN0 ));
 sky130_fd_sc_hd__and3b_2 \BANK128[0].RAM128.DEC0.AND1  (.A_N(\BANK128[0].RAM128.A0BUF[6].X ),
    .B(\BANK128[0].RAM128.A0BUF[5].X ),
    .C(\BANK128[0].RAM128.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[1].RAM32.EN0 ));
 sky130_fd_sc_hd__and3b_2 \BANK128[0].RAM128.DEC0.AND2  (.A_N(\BANK128[0].RAM128.A0BUF[5].X ),
    .B(\BANK128[0].RAM128.A0BUF[6].X ),
    .C(\BANK128[0].RAM128.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[2].RAM32.EN0 ));
 sky130_fd_sc_hd__and3_2 \BANK128[0].RAM128.DEC0.AND3  (.A(\BANK128[0].RAM128.A0BUF[6].X ),
    .B(\BANK128[0].RAM128.A0BUF[5].X ),
    .C(\BANK128[0].RAM128.DEC0.EN ),
    .X(\BANK128[0].RAM128.BLOCK[3].RAM32.EN0 ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.DIBUF[0].__cell__  (.A(Di0[0]),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[0].A ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.DIBUF[1].__cell__  (.A(Di0[1]),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[1].A ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.DIBUF[2].__cell__  (.A(Di0[2]),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[2].A ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.DIBUF[3].__cell__  (.A(Di0[3]),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[3].A ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.DIBUF[4].__cell__  (.A(Di0[4]),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[4].A ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.DIBUF[5].__cell__  (.A(Di0[5]),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[5].A ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.DIBUF[6].__cell__  (.A(Di0[6]),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[6].A ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[0].RAM128.DIBUF[7].__cell__  (.A(Di0[7]),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.DIBUF[7].A ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A0MUX[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A0MUX[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A0MUX[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A0MUX[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A0MUX[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A0MUX[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A0MUX[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A0MUX[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[7] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A1MUX[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A1MUX[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A1MUX[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A1MUX[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A1MUX[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A1MUX[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A1MUX[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A1MUX[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[7] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A2MUX[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A2MUX[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A2MUX[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A2MUX[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A2MUX[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A2MUX[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A2MUX[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A2MUX[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[7] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A3MUX[0]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A3MUX[1]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A3MUX[2]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A3MUX[3]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A3MUX[4]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A3MUX[5]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A3MUX[6]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.M[0].DIODE_A3MUX[7]  (.DIODE(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[7] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[0].RAM128.Do0MUX.M[0].MUX[0]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[0] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[0] ),
    .A2(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[0] ),
    .A3(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[0] ),
    .S0(\BANK128[0].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[0].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[0].RAM128.Do0[0] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[0].RAM128.Do0MUX.M[0].MUX[1]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[1] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[1] ),
    .A2(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[1] ),
    .A3(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[1] ),
    .S0(\BANK128[0].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[0].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[0].RAM128.Do0[1] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[0].RAM128.Do0MUX.M[0].MUX[2]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[2] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[2] ),
    .A2(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[2] ),
    .A3(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[2] ),
    .S0(\BANK128[0].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[0].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[0].RAM128.Do0[2] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[0].RAM128.Do0MUX.M[0].MUX[3]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[3] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[3] ),
    .A2(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[3] ),
    .A3(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[3] ),
    .S0(\BANK128[0].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[0].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[0].RAM128.Do0[3] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[0].RAM128.Do0MUX.M[0].MUX[4]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[4] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[4] ),
    .A2(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[4] ),
    .A3(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[4] ),
    .S0(\BANK128[0].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[0].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[0].RAM128.Do0[4] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[0].RAM128.Do0MUX.M[0].MUX[5]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[5] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[5] ),
    .A2(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[5] ),
    .A3(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[5] ),
    .S0(\BANK128[0].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[0].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[0].RAM128.Do0[5] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[0].RAM128.Do0MUX.M[0].MUX[6]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[6] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[6] ),
    .A2(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[6] ),
    .A3(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[6] ),
    .S0(\BANK128[0].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[0].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[0].RAM128.Do0[6] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[0].RAM128.Do0MUX.M[0].MUX[7]  (.A0(\BANK128[0].RAM128.BLOCK[0].RAM32.Do0[7] ),
    .A1(\BANK128[0].RAM128.BLOCK[1].RAM32.Do0[7] ),
    .A2(\BANK128[0].RAM128.BLOCK[2].RAM32.Do0[7] ),
    .A3(\BANK128[0].RAM128.BLOCK[3].RAM32.Do0[7] ),
    .S0(\BANK128[0].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[0].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[0].RAM128.Do0[7] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.Do0MUX.SEL0BUF[0]  (.A(\BANK128[0].RAM128.A0BUF[5].X ),
    .X(\BANK128[0].RAM128.Do0MUX.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.Do0MUX.SEL1BUF[0]  (.A(\BANK128[0].RAM128.A0BUF[6].X ),
    .X(\BANK128[0].RAM128.Do0MUX.SEL1 ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.SEL_DIODE[0]  (.DIODE(\BANK128[0].RAM128.A0BUF[5].X ));
 sky130_fd_sc_hd__diode_2 \BANK128[0].RAM128.Do0MUX.SEL_DIODE[1]  (.DIODE(\BANK128[0].RAM128.A0BUF[6].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.EN0BUF.__cell__  (.A(\BANK128[0].RAM128.EN0 ),
    .X(\BANK128[0].RAM128.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[0].RAM128.WEBUF[0].__cell__  (.A(WE0),
    .X(\BANK128[0].RAM128.BLOCK[0].RAM32.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.A0BUF[0].__cell__  (.A(A0[0]),
    .X(\BANK128[1].RAM128.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.A0BUF[1].__cell__  (.A(A0[1]),
    .X(\BANK128[1].RAM128.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.A0BUF[2].__cell__  (.A(A0[2]),
    .X(\BANK128[1].RAM128.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.A0BUF[3].__cell__  (.A(A0[3]),
    .X(\BANK128[1].RAM128.A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.A0BUF[4].__cell__  (.A(A0[4]),
    .X(\BANK128[1].RAM128.A0BUF[4].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.A0BUF[5].__cell__  (.A(A0[5]),
    .X(\BANK128[1].RAM128.A0BUF[5].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.A0BUF[6].__cell__  (.A(A0[6]),
    .X(\BANK128[1].RAM128.A0BUF[6].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[0].__cell__  (.A(\BANK128[1].RAM128.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[1].__cell__  (.A(\BANK128[1].RAM128.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[2].__cell__  (.A(\BANK128[1].RAM128.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[3].__cell__  (.A(\BANK128[1].RAM128.A0BUF[3].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[4].__cell__  (.A(\BANK128[1].RAM128.A0BUF[4].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[4].X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.DEC0.AND0  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[4].X ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.EN0 ));
 sky130_fd_sc_hd__and2_2 \BANK128[1].RAM128.BLOCK[0].RAM32.DEC0.AND1  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[4].X ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.EN0 ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].A ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].A ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].A ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].A ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].A ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].A ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].A ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].A ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A0MUX[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].DIODE_A1MUX[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[0]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[0] ),
    .A1(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[0] ),
    .S(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[0] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[1]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[1] ),
    .A1(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[1] ),
    .S(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[1] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[2]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[2] ),
    .A1(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[2] ),
    .S(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[2] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[3]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[3] ),
    .A1(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[3] ),
    .S(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[3] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[4]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[4] ),
    .A1(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[4] ),
    .S(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[4] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[5]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[5] ),
    .A1(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[5] ),
    .S(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[5] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[6]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[6] ),
    .A1(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[6] ),
    .S(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[6] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.M[0].MUX[7]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[7] ),
    .A1(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[7] ),
    .S(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[7] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.SEL0BUF[0]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[4].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.SEL ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.EN0BUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[3].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.DEC0.AND0  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.DEC0.AND1  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.EN0BUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.TIE0[0].__cell__  (.LO(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.A0BUF[3].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.DEC0.AND0  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.DEC0.AND1  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.EN0BUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.TIE0[0].__cell__  (.LO(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[0].RAM32.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.SLICE_16[0].RAM16.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[0].__cell__  (.A(\BANK128[1].RAM128.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[1].__cell__  (.A(\BANK128[1].RAM128.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[2].__cell__  (.A(\BANK128[1].RAM128.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[3].__cell__  (.A(\BANK128[1].RAM128.A0BUF[3].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[4].__cell__  (.A(\BANK128[1].RAM128.A0BUF[4].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[4].X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.DEC0.AND0  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[4].X ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.EN0 ));
 sky130_fd_sc_hd__and2_2 \BANK128[1].RAM128.BLOCK[1].RAM32.DEC0.AND1  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[4].X ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.EN0 ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].A ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].A ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].A ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].A ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].A ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].A ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].A ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].A ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A0MUX[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].DIODE_A1MUX[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[0]  (.A0(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[0] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[0] ),
    .S(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[0] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[1]  (.A0(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[1] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[1] ),
    .S(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[1] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[2]  (.A0(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[2] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[2] ),
    .S(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[2] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[3]  (.A0(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[3] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[3] ),
    .S(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[3] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[4]  (.A0(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[4] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[4] ),
    .S(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[4] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[5]  (.A0(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[5] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[5] ),
    .S(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[5] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[6]  (.A0(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[6] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[6] ),
    .S(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[6] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.M[0].MUX[7]  (.A0(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[7] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[7] ),
    .S(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[7] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.SEL0BUF[0]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[4].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.SEL ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.EN0BUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[3].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.DEC0.AND0  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.DEC0.AND1  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.EN0BUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.TIE0[0].__cell__  (.LO(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.A0BUF[3].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.DEC0.AND0  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.DEC0.AND1  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.EN0BUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.TIE0[0].__cell__  (.LO(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[1].RAM32.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.SLICE_16[0].RAM16.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[0].__cell__  (.A(\BANK128[1].RAM128.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[1].__cell__  (.A(\BANK128[1].RAM128.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[2].__cell__  (.A(\BANK128[1].RAM128.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[3].__cell__  (.A(\BANK128[1].RAM128.A0BUF[3].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[4].__cell__  (.A(\BANK128[1].RAM128.A0BUF[4].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[4].X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.DEC0.AND0  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[4].X ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.EN0 ));
 sky130_fd_sc_hd__and2_2 \BANK128[1].RAM128.BLOCK[2].RAM32.DEC0.AND1  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[4].X ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.EN0 ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].A ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].A ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].A ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].A ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].A ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].A ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].A ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].A ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A0MUX[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].DIODE_A1MUX[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[0]  (.A0(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[0] ),
    .A1(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[0] ),
    .S(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[0] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[1]  (.A0(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[1] ),
    .A1(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[1] ),
    .S(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[1] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[2]  (.A0(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[2] ),
    .A1(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[2] ),
    .S(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[2] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[3]  (.A0(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[3] ),
    .A1(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[3] ),
    .S(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[3] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[4]  (.A0(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[4] ),
    .A1(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[4] ),
    .S(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[4] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[5]  (.A0(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[5] ),
    .A1(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[5] ),
    .S(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[5] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[6]  (.A0(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[6] ),
    .A1(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[6] ),
    .S(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[6] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.M[0].MUX[7]  (.A0(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[7] ),
    .A1(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[7] ),
    .S(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[7] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.SEL0BUF[0]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[4].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.SEL ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.EN0BUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[3].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.DEC0.AND0  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.DEC0.AND1  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.EN0BUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.TIE0[0].__cell__  (.LO(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.A0BUF[3].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.DEC0.AND0  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.DEC0.AND1  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.EN0BUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.TIE0[0].__cell__  (.LO(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[2].RAM32.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.SLICE_16[0].RAM16.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[0].__cell__  (.A(\BANK128[1].RAM128.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[1].__cell__  (.A(\BANK128[1].RAM128.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[2].__cell__  (.A(\BANK128[1].RAM128.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[3].__cell__  (.A(\BANK128[1].RAM128.A0BUF[3].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[4].__cell__  (.A(\BANK128[1].RAM128.A0BUF[4].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[4].X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.DEC0.AND0  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[4].X ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.EN0 ));
 sky130_fd_sc_hd__and2_2 \BANK128[1].RAM128.BLOCK[3].RAM32.DEC0.AND1  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[4].X ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.EN0 ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].A ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].A ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].A ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].A ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].A ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].A ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].A ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].A ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A0MUX[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].DIODE_A1MUX[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[0]  (.A0(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[0] ),
    .A1(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[0] ),
    .S(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[0] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[1]  (.A0(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[1] ),
    .A1(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[1] ),
    .S(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[1] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[2]  (.A0(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[2] ),
    .A1(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[2] ),
    .S(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[2] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[3]  (.A0(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[3] ),
    .A1(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[3] ),
    .S(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[3] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[4]  (.A0(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[4] ),
    .A1(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[4] ),
    .S(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[4] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[5]  (.A0(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[5] ),
    .A1(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[5] ),
    .S(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[5] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[6]  (.A0(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[6] ),
    .A1(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[6] ),
    .S(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[6] ));
 sky130_fd_sc_hd__mux2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.M[0].MUX[7]  (.A0(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[7] ),
    .A1(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[7] ),
    .S(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[7] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.SEL0BUF[0]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[4].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.SEL ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.EN0BUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[3].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.DEC0.AND0  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.DEC0.AND1  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A0[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.EN0BUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.TIE0[0].__cell__  (.LO(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.A0BUF[3].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.CLK ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.CLKBUF.X ));
 sky130_fd_sc_hd__and2b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.DEC0.AND0  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and2_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.DEC0.AND1  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[3].X ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.Do_CLKBUF[0]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLKBUF ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0MUX.A1[7] ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.Root_CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.EN0BUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.FBUFENBUF0[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.EN0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[0].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[1].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.A0BUF[2].X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.AND7  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BANK128[1].RAM128.BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WE0_buf ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.TIE0[0].__cell__  (.LO(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[1].RAM16.SLICE[0].RAM8.WE0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.BLOCK[3].RAM32.WEBUF[0].__cell__  (.A(\BANK128[1].RAM128.BLOCK[0].RAM32.WE0 ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.SLICE_16[0].RAM16.WE0 ));
 sky130_fd_sc_hd__clkbuf_4 \BANK128[1].RAM128.CLKBUF.__cell__  (.A(CLK),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.CLK ));
 sky130_fd_sc_hd__nor3b_2 \BANK128[1].RAM128.DEC0.AND0  (.A(\BANK128[1].RAM128.A0BUF[5].X ),
    .B(\BANK128[1].RAM128.A0BUF[6].X ),
    .C_N(\BANK128[1].RAM128.DEC0.EN ),
    .Y(\BANK128[1].RAM128.BLOCK[0].RAM32.EN0 ));
 sky130_fd_sc_hd__and3b_2 \BANK128[1].RAM128.DEC0.AND1  (.A_N(\BANK128[1].RAM128.A0BUF[6].X ),
    .B(\BANK128[1].RAM128.A0BUF[5].X ),
    .C(\BANK128[1].RAM128.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[1].RAM32.EN0 ));
 sky130_fd_sc_hd__and3b_2 \BANK128[1].RAM128.DEC0.AND2  (.A_N(\BANK128[1].RAM128.A0BUF[5].X ),
    .B(\BANK128[1].RAM128.A0BUF[6].X ),
    .C(\BANK128[1].RAM128.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[2].RAM32.EN0 ));
 sky130_fd_sc_hd__and3_2 \BANK128[1].RAM128.DEC0.AND3  (.A(\BANK128[1].RAM128.A0BUF[6].X ),
    .B(\BANK128[1].RAM128.A0BUF[5].X ),
    .C(\BANK128[1].RAM128.DEC0.EN ),
    .X(\BANK128[1].RAM128.BLOCK[3].RAM32.EN0 ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.DIBUF[0].__cell__  (.A(Di0[0]),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[0].A ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.DIBUF[1].__cell__  (.A(Di0[1]),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[1].A ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.DIBUF[2].__cell__  (.A(Di0[2]),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[2].A ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.DIBUF[3].__cell__  (.A(Di0[3]),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[3].A ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.DIBUF[4].__cell__  (.A(Di0[4]),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[4].A ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.DIBUF[5].__cell__  (.A(Di0[5]),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[5].A ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.DIBUF[6].__cell__  (.A(Di0[6]),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[6].A ));
 sky130_fd_sc_hd__clkbuf_16 \BANK128[1].RAM128.DIBUF[7].__cell__  (.A(Di0[7]),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.DIBUF[7].A ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A0MUX[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A0MUX[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A0MUX[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A0MUX[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A0MUX[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A0MUX[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A0MUX[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A0MUX[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[7] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A1MUX[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A1MUX[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A1MUX[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A1MUX[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A1MUX[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A1MUX[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A1MUX[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A1MUX[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[7] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A2MUX[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A2MUX[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A2MUX[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A2MUX[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A2MUX[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A2MUX[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A2MUX[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A2MUX[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[7] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A3MUX[0]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[0] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A3MUX[1]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[1] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A3MUX[2]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[2] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A3MUX[3]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[3] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A3MUX[4]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[4] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A3MUX[5]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[5] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A3MUX[6]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[6] ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.M[0].DIODE_A3MUX[7]  (.DIODE(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[7] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[1].RAM128.Do0MUX.M[0].MUX[0]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[0] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[0] ),
    .A2(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[0] ),
    .A3(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[0] ),
    .S0(\BANK128[1].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[1].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[1].RAM128.Do0[0] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[1].RAM128.Do0MUX.M[0].MUX[1]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[1] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[1] ),
    .A2(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[1] ),
    .A3(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[1] ),
    .S0(\BANK128[1].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[1].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[1].RAM128.Do0[1] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[1].RAM128.Do0MUX.M[0].MUX[2]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[2] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[2] ),
    .A2(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[2] ),
    .A3(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[2] ),
    .S0(\BANK128[1].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[1].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[1].RAM128.Do0[2] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[1].RAM128.Do0MUX.M[0].MUX[3]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[3] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[3] ),
    .A2(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[3] ),
    .A3(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[3] ),
    .S0(\BANK128[1].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[1].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[1].RAM128.Do0[3] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[1].RAM128.Do0MUX.M[0].MUX[4]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[4] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[4] ),
    .A2(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[4] ),
    .A3(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[4] ),
    .S0(\BANK128[1].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[1].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[1].RAM128.Do0[4] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[1].RAM128.Do0MUX.M[0].MUX[5]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[5] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[5] ),
    .A2(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[5] ),
    .A3(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[5] ),
    .S0(\BANK128[1].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[1].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[1].RAM128.Do0[5] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[1].RAM128.Do0MUX.M[0].MUX[6]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[6] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[6] ),
    .A2(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[6] ),
    .A3(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[6] ),
    .S0(\BANK128[1].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[1].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[1].RAM128.Do0[6] ));
 sky130_fd_sc_hd__mux4_1 \BANK128[1].RAM128.Do0MUX.M[0].MUX[7]  (.A0(\BANK128[1].RAM128.BLOCK[0].RAM32.Do0[7] ),
    .A1(\BANK128[1].RAM128.BLOCK[1].RAM32.Do0[7] ),
    .A2(\BANK128[1].RAM128.BLOCK[2].RAM32.Do0[7] ),
    .A3(\BANK128[1].RAM128.BLOCK[3].RAM32.Do0[7] ),
    .S0(\BANK128[1].RAM128.Do0MUX.SEL0 ),
    .S1(\BANK128[1].RAM128.Do0MUX.SEL1 ),
    .X(\BANK128[1].RAM128.Do0[7] ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.Do0MUX.SEL0BUF[0]  (.A(\BANK128[1].RAM128.A0BUF[5].X ),
    .X(\BANK128[1].RAM128.Do0MUX.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.Do0MUX.SEL1BUF[0]  (.A(\BANK128[1].RAM128.A0BUF[6].X ),
    .X(\BANK128[1].RAM128.Do0MUX.SEL1 ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.SEL_DIODE[0]  (.DIODE(\BANK128[1].RAM128.A0BUF[5].X ));
 sky130_fd_sc_hd__diode_2 \BANK128[1].RAM128.Do0MUX.SEL_DIODE[1]  (.DIODE(\BANK128[1].RAM128.A0BUF[6].X ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.EN0BUF.__cell__  (.A(\BANK128[1].RAM128.EN0 ),
    .X(\BANK128[1].RAM128.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BANK128[1].RAM128.WEBUF[0].__cell__  (.A(WE0),
    .X(\BANK128[1].RAM128.BLOCK[0].RAM32.WE0 ));
 sky130_fd_sc_hd__and2b_2 \DEC0.AND0  (.A_N(A0[7]),
    .B(EN0),
    .X(\BANK128[0].RAM128.EN0 ));
 sky130_fd_sc_hd__and2_2 \DEC0.AND1  (.A(A0[7]),
    .B(EN0),
    .X(\BANK128[1].RAM128.EN0 ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[0]  (.DIODE(\BANK128[0].RAM128.Do0[0] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[1]  (.DIODE(\BANK128[0].RAM128.Do0[1] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[2]  (.DIODE(\BANK128[0].RAM128.Do0[2] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[3]  (.DIODE(\BANK128[0].RAM128.Do0[3] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[4]  (.DIODE(\BANK128[0].RAM128.Do0[4] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[5]  (.DIODE(\BANK128[0].RAM128.Do0[5] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[6]  (.DIODE(\BANK128[0].RAM128.Do0[6] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[7]  (.DIODE(\BANK128[0].RAM128.Do0[7] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[0]  (.DIODE(\BANK128[1].RAM128.Do0[0] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[1]  (.DIODE(\BANK128[1].RAM128.Do0[1] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[2]  (.DIODE(\BANK128[1].RAM128.Do0[2] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[3]  (.DIODE(\BANK128[1].RAM128.Do0[3] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[4]  (.DIODE(\BANK128[1].RAM128.Do0[4] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[5]  (.DIODE(\BANK128[1].RAM128.Do0[5] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[6]  (.DIODE(\BANK128[1].RAM128.Do0[6] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[7]  (.DIODE(\BANK128[1].RAM128.Do0[7] ));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[0]  (.A0(\BANK128[0].RAM128.Do0[0] ),
    .A1(\BANK128[1].RAM128.Do0[0] ),
    .S(\Do0MUX.SEL ),
    .X(Do0[0]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[1]  (.A0(\BANK128[0].RAM128.Do0[1] ),
    .A1(\BANK128[1].RAM128.Do0[1] ),
    .S(\Do0MUX.SEL ),
    .X(Do0[1]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[2]  (.A0(\BANK128[0].RAM128.Do0[2] ),
    .A1(\BANK128[1].RAM128.Do0[2] ),
    .S(\Do0MUX.SEL ),
    .X(Do0[2]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[3]  (.A0(\BANK128[0].RAM128.Do0[3] ),
    .A1(\BANK128[1].RAM128.Do0[3] ),
    .S(\Do0MUX.SEL ),
    .X(Do0[3]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[4]  (.A0(\BANK128[0].RAM128.Do0[4] ),
    .A1(\BANK128[1].RAM128.Do0[4] ),
    .S(\Do0MUX.SEL ),
    .X(Do0[4]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[5]  (.A0(\BANK128[0].RAM128.Do0[5] ),
    .A1(\BANK128[1].RAM128.Do0[5] ),
    .S(\Do0MUX.SEL ),
    .X(Do0[5]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[6]  (.A0(\BANK128[0].RAM128.Do0[6] ),
    .A1(\BANK128[1].RAM128.Do0[6] ),
    .S(\Do0MUX.SEL ),
    .X(Do0[6]));
 sky130_fd_sc_hd__mux2_1 \Do0MUX.M[0].MUX[7]  (.A0(\BANK128[0].RAM128.Do0[7] ),
    .A1(\BANK128[1].RAM128.Do0[7] ),
    .S(\Do0MUX.SEL ),
    .X(Do0[7]));
 sky130_fd_sc_hd__clkbuf_2 \Do0MUX.SEL0BUF[0]  (.A(A0[7]),
    .X(\Do0MUX.SEL ));

endmodule

