// tb_carry_lookahead_toplayici.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module tb_carry_lookahead_toplayici();

    carry_lookahead_toplayici clat(

    );

    initial begin

        $finish;
    end

endmodule
