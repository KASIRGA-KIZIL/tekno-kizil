// tb_sifreleme_birimi.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module tb_sifreleme_birimi();

    sifreleme_birimi sb(

    );

    initial begin

        $finish;
    end

endmodule
