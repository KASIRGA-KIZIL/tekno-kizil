// OpenRAM SRAM model
// Words: 512
// Word size: 41

module sram_41_512_sky130(
`ifdef USE_POWER_PINS
    vccd1,
    vssd1,
`endif
// Port 0: W
    clk0,csb0,spare_wen0,addr0,din0,
// Port 1: // OpenRAM SRAM model
// Words: 512
// Word size: 54

module sram_54b_512_1w_1r_sky130(
  `ifdef USE_POWER_PINS
      vccd1,
      vssd1,
  `endif
  // Port 0: W
      clk0,csb0,spare_wen0,addr0,din0,
  // Port 1: R
      clk1,csb1,addr1,dout1
    );
  
    parameter DATA_WIDTH = 55 ;
    parameter ADDR_WIDTH = 9 ;
    parameter RAM_DEPTH = 1 << ADDR_WIDTH;
    // FIXME: This delay is arbitrary.
    parameter DELAY = 3 ;
    parameter VERBOSE = 1 ; //Set to 0 to only display warnings
    parameter T_HOLD = 1 ; //Delay to hold dout value after posedge. Value is arbitrary
  
  `ifdef USE_POWER_PINS
      inout vccd1;
      inout vssd1;
  `endif
    input  clk0; // clock
    input   csb0; // active low chip select
    input [ADDR_WIDTH-1:0]  addr0;
    input           spare_wen0; // spare mask
    input [DATA_WIDTH-1:0]  din0;
    input  clk1; // clock
    input   csb1; // active low chip select
    input [ADDR_WIDTH-1:0]  addr1;
    output [DATA_WIDTH-1:0] dout1;
  
    reg [DATA_WIDTH-1:0]    mem [0:RAM_DEPTH-1];
  
    reg  csb0_reg;
    reg spare_wen0_reg;
    reg [ADDR_WIDTH-1:0]  addr0_reg;
    reg [DATA_WIDTH-1:0]  din0_reg;
  
    // All inputs are registers
    always @(posedge clk0)
    begin
      csb0_reg = csb0;
      spare_wen0_reg = spare_wen0;
      addr0_reg = addr0;
      din0_reg = din0;
      if ( !csb0_reg && VERBOSE )
        $display($time," Writing %m addr0=%b din0=%b",addr0_reg,din0_reg);
    end
  
    reg  csb1_reg;
    reg [ADDR_WIDTH-1:0]  addr1_reg;
    reg [DATA_WIDTH-1:0]  dout1;
  
    // All inputs are registers
    always @(posedge clk1)
    begin
      csb1_reg = csb1;
      addr1_reg = addr1;
      if (!csb0 && !csb1 && (addr0 == addr1))
           $display($time," WARNING: Writing and reading addr0=%b and addr1=%b simultaneously!",addr0,addr1);
      #(T_HOLD) dout1 = 54'bx;
      if ( !csb1_reg && VERBOSE ) 
        $display($time," Reading %m addr1=%b dout1=%b",addr1_reg,mem[addr1_reg]);
    end
  
  
    // Memory Write Block Port 0
    // Write Operation : When web0 = 0, csb0 = 0
    always @ (negedge clk0)
    begin : MEM_WRITE0
      if (!csb0_reg) begin
          mem[addr0_reg][52:0] = din0_reg[52:0];
          if (spare_wen0_reg)
                  mem[addr0_reg][54] = din0_reg[54];
      end
    end
  
    // Memory Read Block Port 1
    // Read Operation : When web1 = 1, csb1 = 0
    always @ (negedge clk1)
    begin : MEM_READ1
      if (!csb1_reg)
         dout1 <= #(DELAY) mem[addr1_reg];
    end
  
  endmodule
    clk1,csb1,addr1,dout1
  );

  parameter DATA_WIDTH = 42 ;
  parameter ADDR_WIDTH = 9 ;
  parameter RAM_DEPTH = 1 << ADDR_WIDTH;
  // FIXME: This delay is arbitrary.
  parameter DELAY = 3 ;
  parameter VERBOSE = 0 ; //Set to 0 to only display warnings
  parameter T_HOLD = 1 ; //Delay to hold dout value after posedge. Value is arbitrary

`ifdef USE_POWER_PINS
    inout vccd1;
    inout vssd1;
`endif
  input  clk0; // clock
  input   csb0; // active low chip select
  input [ADDR_WIDTH-1:0]  addr0;
  input           spare_wen0; // spare mask
  input [DATA_WIDTH-1:0]  din0;
  input  clk1; // clock
  input   csb1; // active low chip select
  input [ADDR_WIDTH-1:0]  addr1;
  output [DATA_WIDTH-1:0] dout1;

  reg [DATA_WIDTH-1:0]    mem [0:RAM_DEPTH-1];

  reg  csb0_reg;
  reg spare_wen0_reg;
  reg [ADDR_WIDTH-1:0]  addr0_reg;
  reg [DATA_WIDTH-1:0]  din0_reg;

  // All inputs are registers
  always @(posedge clk0)
  begin
    csb0_reg = csb0;
    spare_wen0_reg = spare_wen0;
    addr0_reg = addr0;
    din0_reg = din0;
    if ( !csb0_reg && VERBOSE )
      $display($time," Writing %m addr0=%b din0=%b",addr0_reg,din0_reg);
  end

  reg  csb1_reg;
  reg [ADDR_WIDTH-1:0]  addr1_reg;
  reg [DATA_WIDTH-1:0]  dout1;

  // All inputs are registers
  always @(posedge clk1)
  begin
    csb1_reg = csb1;
    addr1_reg = addr1;
    if (!csb0 && !csb1 && (addr0 == addr1))
         $display($time," WARNING: Writing and reading addr0=%b and addr1=%b simultaneously!",addr0,addr1);
    #(T_HOLD) dout1 = 41'bx;
    if ( !csb1_reg && VERBOSE )
      $display($time," Reading %m addr1=%b dout1=%b",addr1_reg,mem[addr1_reg]);
  end


  // Memory Write Block Port 0
  // Write Operation : When web0 = 0, csb0 = 0
  always @ (negedge clk0)
  begin : MEM_WRITE0
    if (!csb0_reg) begin
        mem[addr0_reg][39:0] = din0_reg[39:0];
        if (spare_wen0_reg)
                mem[addr0_reg][41] = din0_reg[41];
    end
  end

  // Memory Read Block Port 1
  // Read Operation : When web1 = 1, csb1 = 0
  always @ (negedge clk1)
  begin : MEM_READ1
    if (!csb1_reg)
       dout1 <= #(DELAY) mem[addr1_reg];
  end

endmodule
