// tb_modified_booth_dadda_carpici.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module tb_modified_booth_dadda_carpici();

    modified_booth_dadda_carpici mbdc(

    );

    initial begin

        $finish;
    end

endmodule
