@40000000
13 01 01 FF 23 26 11 00 23 24 81 00 EF 00 50 3C
17 15 00 00 13 05 45 C0 EF 00 C0 2D 17 15 00 00
13 05 05 C0 EF 00 00 2D EF 00 10 3D EF 00 D0 3C
EF 00 90 3C EF 00 50 3C 17 15 00 00 13 05 C5 BE
EF 00 40 2B 17 14 00 00 13 04 44 BE EF 00 D0 3A
93 05 05 00 13 05 04 00 EF 00 C0 29 6F F0 1F FF
6F 00 00 00 13 01 01 FA 23 2E 81 04 23 2C 91 04
13 F8 07 04 97 1E 00 00 93 8E 0E BE 63 16 08 00
97 1E 00 00 93 8E CE BA 13 F4 07 01 63 16 04 14
13 F8 17 00 93 F4 17 01 93 03 00 03 63 02 08 14
13 F8 27 00 13 FF 07 02 63 04 08 12 63 C4 05 14
13 F8 47 00 63 14 08 18 93 F7 87 00 93 0F 00 00
63 86 07 00 93 86 F6 FF 93 0F 00 02 63 0C 0F 00
93 07 00 01 63 0E F6 18 93 07 86 FF 93 B7 17 00
B3 86 F6 40 63 90 05 12 93 07 00 03 23 06 F1 00
13 08 10 00 93 02 C1 00 93 08 08 00 63 54 E8 00
93 08 07 00 B3 86 16 41 63 90 04 02 33 07 D5 00
93 07 00 02 63 5A D0 16 13 05 15 00 A3 0F F5 FE
E3 1C E5 FE 93 06 F0 FF 63 86 0F 00 23 00 F5 01
13 05 15 00 63 0A 0F 00 93 07 80 00 63 02 F6 12
93 07 00 01 63 02 F6 10 63 1E 04 00 B3 07 D5 00
63 50 D0 14 13 05 15 00 A3 0F 75 FE E3 9C A7 FE
93 06 F0 FF B3 87 08 41 B3 07 F5 00 13 07 00 03
63 58 18 11 13 05 15 00 A3 0F E5 FE E3 9C A7 FE
33 87 B2 00 13 86 07 00 03 48 07 00 13 05 07 00
13 06 16 00 A3 0F 06 FF 13 07 F7 FF E3 96 A2 FE
93 85 15 00 B3 85 B7 00 63 58 D0 0C 33 85 D5 00
93 07 00 02 93 85 15 00 A3 8F F5 FE E3 1C B5 FE
03 24 C1 05 83 24 81 05 13 01 01 06 67 80 00 00
93 0F 00 00 6F F0 9F EF 93 F7 E7 FF 93 04 04 00
13 F8 27 00 93 03 00 02 13 FF 07 02 E3 02 08 FE
6F F0 DF EB B3 05 B0 40 93 86 F6 FF 93 0F D0 02
E3 18 0F EC 93 87 05 00 13 08 00 00 93 02 C1 00
B3 F8 C7 02 93 05 08 00 13 08 18 00 33 8E 02 01
13 83 07 00 B3 88 1E 01 83 C8 08 00 B3 D7 C7 02
A3 0F 1E FF E3 7E C3 FC 6F F0 1F EC 93 86 F6 FF
93 0F B0 02 6F F0 9F E8 93 07 00 03 23 00 F5 00
93 07 80 07 A3 00 F5 00 13 05 25 00 6F F0 DF EE
93 07 00 03 23 00 F5 00 13 05 15 00 6F F0 DF ED
93 86 E6 FF 6F F0 1F E7 13 85 05 00 6F F0 5F F4
93 07 05 00 6F F0 DF EF 93 86 F6 FF 6F F0 DF E9
93 86 F6 FF 6F F0 1F ED 37 07 00 20 83 27 47 00
93 F7 17 00 E3 9C 07 FE 23 06 A7 00 67 80 00 00
83 46 05 00 63 82 06 02 37 07 00 20 13 05 15 00
83 27 47 00 93 F7 17 00 E3 9C 07 FE 23 06 D7 00
83 46 05 00 E3 94 06 FE 67 80 00 00 37 07 00 20
83 27 47 00 93 F7 17 00 E3 9C 07 FE 23 06 A7 00
67 80 00 00 13 01 01 B7 23 20 E1 48 23 26 11 46
23 24 81 46 23 22 91 46 23 20 21 47 23 2E 31 45
23 2C 41 45 23 2A 51 45 23 28 61 45 23 26 71 45
23 24 81 45 23 22 91 45 23 20 A1 45 23 2E B1 43
23 2A B1 46 23 2C C1 46 23 2E D1 46 23 22 F1 48
23 24 01 49 23 26 11 49 83 47 05 00 13 07 41 47
23 2A E1 00 63 8A 07 72 93 09 01 03 13 03 05 00
13 0A 07 00 13 85 09 00 13 09 50 02 93 04 00 01
17 14 00 00 13 04 44 91 93 0D 90 00 93 0C E0 02
13 0D C0 04 13 0C 70 03 63 88 27 05 23 00 F5 00
83 47 13 00 13 05 15 00 13 03 13 00 E3 96 07 FE
23 00 05 00 03 46 01 03 63 08 06 10 93 86 09 00
37 07 00 20 83 27 47 00 93 F7 17 00 E3 9C 07 FE
23 06 C7 00 03 C6 16 00 93 87 16 00 63 04 06 12
93 86 07 00 6F F0 1F FE 93 07 00 00 03 46 13 00
93 05 13 00 13 07 06 FE 13 77 F7 0F 63 EC E4 00
13 17 27 00 33 07 87 00 03 27 07 00 33 07 87 00
67 00 07 00 13 07 06 FD 13 77 F7 0F 63 FC ED 14
13 07 A0 02 93 06 F0 FF 63 00 E6 18 13 07 F0 FF
63 0C 96 11 13 78 F6 0D 63 0C A8 09 13 08 F6 FB
13 78 F8 0F 63 6E 0C 05 97 18 00 00 93 88 08 89
13 18 28 00 33 08 18 01 03 28 08 00 33 08 18 01
67 00 08 00 93 E7 17 00 13 83 05 00 6F F0 1F F8
93 E7 07 01 13 83 05 00 6F F0 5F F7 93 E7 47 00
13 83 05 00 6F F0 9F F6 93 E7 07 02 13 83 05 00
6F F0 DF F5 93 E7 87 00 13 83 05 00 6F F0 1F F5
93 8A 05 00 93 07 50 02 63 04 F6 58 23 00 F5 00
83 C7 0A 00 13 05 15 00 63 9E 07 56 23 00 05 00
03 46 01 03 E3 1C 06 EE 13 05 00 00 6F 00 00 04
93 08 06 00 03 C6 15 00 93 8A 15 00 13 08 F6 FB
13 78 F8 0F E3 60 0C FD 17 13 00 00 13 03 03 8D
13 18 28 00 33 08 68 00 03 28 08 00 33 08 68 00
67 00 08 00 B3 86 36 41 13 85 16 00 83 20 C1 46
03 24 81 46 83 24 41 46 03 29 01 46 83 29 C1 45
03 2A 81 45 83 2A 41 45 03 2B 01 45 83 2B C1 44
03 2C 81 44 83 2C 41 44 03 2D 01 44 83 2D C1 43
13 01 01 49 67 80 00 00 03 C6 15 00 93 08 90 00
13 88 15 00 13 07 06 FD 13 77 F7 0F 63 FA E8 36
13 07 A0 02 63 04 E6 3A 93 05 08 00 13 07 00 00
6F F0 5F EC 93 06 00 00 13 08 90 00 13 97 26 00
33 07 D7 00 93 85 15 00 13 17 17 00 33 07 C7 00
03 C6 05 00 93 06 07 FD 13 07 06 FD 13 77 F7 0F
E3 7E E8 FC 6F F0 9F E8 83 26 0A 00 03 46 23 00
93 05 23 00 13 0A 4A 00 E3 DA 06 E6 B3 06 D0 40
93 E7 07 01 6F F0 9F E6 93 E7 07 04 13 07 C0 06
63 80 E8 36 03 2E 0A 00 93 05 00 00 13 07 00 00
33 06 BE 00 03 46 06 00 23 24 F1 00 23 26 D1 00
93 0F 4A 00 93 03 30 06 97 0E 00 00 93 8E 4E 64
13 0B 40 06 93 0B A0 00 93 02 00 03 13 03 40 00
13 0F E0 02 13 08 17 00 63 10 06 04 93 07 07 42
13 07 01 01 33 87 E7 00 23 04 57 BE 93 85 15 00
63 82 65 0A 93 07 08 42 13 07 01 01 33 86 E7 00
23 04 E6 BF 33 06 BE 00 03 46 06 00 13 07 18 00
13 08 17 00 E3 04 06 FC 63 DA C3 22 B3 67 66 03
93 06 07 42 93 08 01 01 B3 88 16 01 93 86 08 00
13 08 08 42 93 08 01 01 33 08 18 01 23 22 01 01
13 07 27 00 93 88 0E 00 13 08 17 00 33 46 66 03
33 CA 77 03 33 86 CE 00 03 46 06 00 23 84 C6 BE
33 8A 4E 01 33 E6 77 03 03 4A 0A 00 83 27 41 00
23 84 47 BF B3 88 C8 00 03 C6 08 00 93 07 07 42
13 07 01 01 33 87 E7 00 23 04 C7 BE 93 85 15 00
E3 92 65 F6 83 27 81 00 83 26 C1 00 93 F7 07 01
63 96 07 02 13 86 F6 FF 63 5E D8 4A B3 87 06 41
B3 07 F5 00 13 07 00 02 13 05 15 00 A3 0F E5 FE
E3 9C A7 FE B3 06 D8 40 B3 86 C6 00 13 06 81 01
B3 07 05 01 13 07 05 00 83 45 06 00 13 07 17 00
13 06 16 00 A3 0F B7 FE E3 98 E7 FE 63 58 D8 44
33 05 D5 00 13 07 00 02 93 87 17 00 A3 8F E7 FE
E3 9C A7 FE 83 C7 1A 00 13 83 1A 00 13 8A 0F 00
E3 94 07 C4 6F F0 DF C5 93 E7 07 04 13 06 00 01
13 08 4A 00 83 25 0A 00 13 0A 08 00 EF F0 9F 90
83 C7 1A 00 13 83 1A 00 E3 90 07 C2 6F F0 5F C3
93 8A 05 00 93 F7 07 01 13 06 4A 00 13 83 1A 00
63 8A 07 2C 83 27 0A 00 93 05 10 00 13 07 15 00
23 00 F5 00 93 07 00 02 33 05 D5 00 63 D4 D5 40
13 07 17 00 A3 0F F7 FE E3 1C A7 FE 83 C7 1A 00
13 0A 06 00 E3 9A 07 BC 6F F0 9F BE 93 8A 05 00
03 26 0A 00 13 0A 4A 00 63 00 06 28 83 45 06 00
63 8E 05 30 63 0C 07 30 93 05 06 00 6F 00 C0 00
33 88 E5 40 63 08 C8 00 03 C8 15 00 93 85 15 00
E3 18 08 FE 13 F7 07 01 B3 87 C5 40 63 0C 07 28
63 5C F0 3A 33 08 F6 00 13 07 05 00 83 45 06 00
13 06 16 00 13 07 17 00 A3 0F B7 FE E3 18 06 FF
33 07 F5 00 33 85 F6 40 13 83 1A 00 33 05 A7 00
13 06 00 02 63 D8 D7 34 13 07 17 00 A3 0F C7 FE
E3 1C A7 FE 83 C7 1A 00 E3 90 07 B4 6F F0 5F B5
93 8A 05 00 13 06 F0 FF 63 82 C6 1E 83 25 0A 00
13 06 00 01 13 0A 4A 00 EF F0 CF FF 83 C7 1A 00
13 83 1A 00 E3 9A 07 B0 6F F0 9F B2 93 07 90 00
93 88 0E 00 E3 D0 C7 E2 13 0A A0 00 B3 47 46 03
97 08 00 00 93 88 C8 39 13 07 07 42 93 06 01 01
B3 06 D7 00 13 07 08 00 13 08 18 00 33 66 46 03
33 8A F8 00 03 4A 0A 00 23 84 46 BF 6F F0 9F DE
13 07 00 00 13 03 07 00 13 17 23 00 33 07 67 00
13 08 18 00 13 17 17 00 33 07 C7 00 03 46 08 00
13 03 07 FD 93 05 06 FD 93 F5 F5 0F E3 FE B8 FC
13 07 03 00 93 05 08 00 6F F0 DF B2 03 27 0A 00
13 88 25 00 03 C6 25 00 93 45 F7 FF 93 D5 F5 41
33 77 B7 00 13 0A 4A 00 93 05 08 00 6F F0 9F B0
13 F7 07 04 17 03 00 00 13 03 83 30 63 06 07 00
17 03 00 00 13 03 43 32 83 2E 0A 00 13 06 00 00
93 08 00 00 13 0E 60 00 13 0F A0 03 6F 00 40 01
13 87 28 42 33 08 77 00 93 88 38 00 23 04 E8 BF
33 87 CE 00 03 47 07 00 93 03 01 01 13 06 16 00
13 58 47 00 13 77 F7 00 33 07 E3 00 33 08 03 01
83 4F 07 00 83 42 08 00 13 87 08 42 33 07 77 00
23 04 57 BE A3 04 F7 BF E3 1C C6 FB 93 F7 07 01
63 98 07 02 93 07 10 01 13 86 F6 FF 63 DE D7 20
93 87 F6 FE B3 07 F5 00 13 07 00 02 13 05 15 00
A3 0F E5 FE E3 9C A7 FE 33 06 D6 40 93 06 16 01
13 06 81 01 93 07 15 01 13 07 05 00 03 48 06 00
13 07 17 00 13 06 16 00 A3 0F 07 FF E3 18 F7 FE
13 06 10 01 63 54 D6 1A 33 05 D5 00 13 07 00 02
93 87 17 00 A3 8F E7 FE E3 1C F5 FE 83 C7 25 00
13 0A 4A 00 13 83 25 00 E3 98 07 96 6F F0 5F 98
83 C7 0A 00 23 00 F5 00 83 C7 1A 00 13 05 15 00
13 83 1A 00 E3 9A 07 94 6F F0 9F 96 93 E7 17 00
93 06 80 00 6F F0 9F E1 17 06 00 00 13 06 46 23
6F F0 5F D8 93 07 10 00 63 DC D7 0E 93 87 F6 FF
B3 07 F5 00 13 07 00 02 13 05 15 00 A3 0F E5 FE
E3 1C F5 FE 93 06 00 00 6F F0 DF D0 93 E7 27 00
13 06 A0 00 6F F0 DF CC 93 09 01 03 13 85 09 00
6F F0 1F 91 13 88 F6 FF 63 D4 D7 12 33 87 F6 40
33 07 E5 00 93 05 00 02 13 05 15 00 A3 0F B5 FE
E3 1C E5 FE B3 86 D7 40 B3 86 06 01 6F F0 5F D4
93 E7 27 00 13 08 4A 00 93 8A 05 00 13 06 A0 00
6F F0 5F C8 13 06 80 00 6F F0 9F C7 13 06 A0 00
6F F0 1F C7 93 8A 05 00 6F F0 DF AD 93 F7 07 01
63 82 07 08 13 07 05 00 93 07 00 00 6F F0 9F D2
93 E7 07 04 93 8A 05 00 6F F0 DF AB 13 08 4A 00
93 8A 05 00 13 06 A0 00 6F F0 DF C3 93 E7 07 04
13 08 4A 00 93 8A 05 00 13 06 00 01 6F F0 9F C2
13 08 4A 00 93 8A 05 00 13 06 00 01 6F F0 9F C1
13 08 4A 00 93 8A 05 00 13 06 80 00 6F F0 9F C0
83 27 0A 00 13 05 15 00 13 0A 06 00 A3 0F F5 FE
83 C7 1A 00 E3 92 07 82 6F F0 9F 83 13 85 07 00
6F F0 5F BC 13 88 F6 FF E3 42 D0 F2 13 83 1A 00
13 07 05 00 83 C7 1A 00 13 05 07 00 63 9E 07 FE
6F F0 1F 81 93 06 06 00 6F F0 5F B6 13 05 07 00
6F F0 DF E6 83 C7 1A 00 13 0A 06 00 13 05 07 00
63 9C 07 FC 6F F0 CF FE 13 07 05 00 6F F0 9F C6
93 06 08 00 6F F0 DF C3 93 06 06 00 6F F0 5F E0
B7 07 00 20 03 A7 07 00 13 67 17 00 23 A0 E7 00
03 A7 07 00 13 67 27 00 23 A0 E7 00 13 07 D0 43
23 91 E7 00 67 80 00 00 37 07 00 20 83 27 47 00
93 D7 37 00 93 F7 17 00 E3 9A 07 FE 03 45 87 00
67 80 00 00
@40000C14
68 65 6C 6C 6F 00 00 00 64 6F 6E 65 00 00 00 00
66 00 00 00 25 63 00 00 30 31 32 33 34 35 36 37
38 39 61 62 63 64 65 66 67 68 69 6A 6B 6C 6D 6E
6F 70 71 72 73 74 75 76 77 78 79 7A 00 00 00 00
30 31 32 33 34 35 36 37 38 39 41 42 43 44 45 46
47 48 49 4A 4B 4C 4D 4E 4F 50 51 52 53 54 55 56
57 58 59 5A 00 00 00 00 3C 4E 55 4C 4C 3E 00
@40000C84
00 F8 FF FF 80 F7 FF FF 80 F7 FF FF F4 F7 FF FF
80 F7 FF FF 80 F7 FF FF 80 F7 FF FF 80 F7 FF FF
80 F7 FF FF 80 F7 FF FF 80 F7 FF FF E8 F7 FF FF
80 F7 FF FF DC F7 FF FF 80 F7 FF FF 80 F7 FF FF
D0 F7 FF FF 38 FE FF FF C8 F7 FF FF C8 F7 FF FF
C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF
C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF
C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF
C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF
C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF
54 FE FF FF C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF
C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF
C8 F7 FF FF 1C FE FF FF C8 F7 FF FF A8 FA FF FF
F8 FD FF FF C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF
C8 F7 FF FF F8 FD FF FF C8 F7 FF FF C8 F7 FF FF
C8 F7 FF FF C8 F7 FF FF C8 F7 FF FF 78 FE FF FF
88 FB FF FF C8 F7 FF FF C8 F7 FF FF F4 FA FF FF
C8 F7 FF FF 44 FE FF FF C8 F7 FF FF C8 F7 FF FF
68 FE FF FF 10 F8 FF FF EC F6 FF FF EC F6 FF FF
EC F6 FF FF EC F6 FF FF EC F6 FF FF EC F6 FF FF
EC F6 FF FF EC F6 FF FF EC F6 FF FF EC F6 FF FF
EC F6 FF FF EC F6 FF FF EC F6 FF FF EC F6 FF FF
EC F6 FF FF EC F6 FF FF EC F6 FF FF EC F6 FF FF
EC F6 FF FF EC F6 FF FF EC F6 FF FF EC F6 FF FF
A0 F9 FF FF EC F6 FF FF EC F6 FF FF EC F6 FF FF
EC F6 FF FF EC F6 FF FF EC F6 FF FF EC F6 FF FF
EC F6 FF FF 14 F8 FF FF EC F6 FF FF CC F9 FF FF
D4 FC FF FF EC F6 FF FF EC F6 FF FF EC F6 FF FF
EC F6 FF FF D4 FC FF FF EC F6 FF FF EC F6 FF FF
EC F6 FF FF EC F6 FF FF EC F6 FF FF 2C FD FF FF
AC FA FF FF EC F6 FF FF EC F6 FF FF 18 FA FF FF
EC F6 FF FF 34 FD FF FF EC F6 FF FF EC F6 FF FF
A4 F9 FF FF
