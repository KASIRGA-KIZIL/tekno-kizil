// aritmetik_mantik_birimi.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module aritmetik_mantik_birimi(


);


endmodule
