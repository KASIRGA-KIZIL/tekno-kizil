// yazmacoku_yurut.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module yazmacoku_yurut(
    input clk_i,
    input rst_i


);


endmodule
