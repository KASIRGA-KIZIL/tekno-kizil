// Toplam 87 buyruk

`define GECERSIZ 7'b0000000

`define ADD_MI 7'b0000010
`define ADDI_MI 7'b0000011
`define AND_MI 7'b0000100
`define ANDI_MI 7'b0000101
`define AUIPC_MI 7'b0000110
`define BEQ_MI 7'b0000111
`define BGE_MI 7'b0001000
`define BGEU_MI 7'b0001001
`define BLT_MI 7'b0001010
`define BLTU_MI 7'b0001011
`define BNE_MI 7'b0001100

`define C_ADD_MI 7'b0001101
`define C_ADDI_MI 7'b0001110
`define C_ADDI16SP_MI 7'b0001111
`define C_ADDI4SPN_MI 7'b0010000
`define C_AND_MI 7'b0010001
`define C_ANDI_MI 7'b0010010
`define C_BEQZ_MI 7'b0010011
`define C_BNEZ_MI 7'b0010100
`define C_EBREAK_MI 7'b0010101
`define C_J_MI 7'b0010110
`define C_JAL_MI 7'b0010111
`define C_JALR_MI 7'b0011000
`define C_JR_MI 7'b0011001
`define C_LI_MI 7'b0011010
`define C_LUI_MI 7'b0011011
`define C_LW_MI 7'b0011100
`define C_LWSP_MI 7'b0011101
`define C_MV_MI 7'b0011110
`define C_NOP_MI 7'b0011111
`define C_OR_MI 7'b0100000
`define C_SLLI_MI 7'b0100001
`define C_SRAI_MI 7'b0100010
`define C_SRLI_MI 7'b0100011
`define C_SUB_MI 7'b0100100
`define C_SW_MI 7'b0100101
`define C_SWSP_MI 7'b0100110
`define C_XOR_MI 7'b0100111

`define DIV_MI 7'b0101000
`define DIVU_MI 7'b0101001
`define EBREAK_MI 7'b0101010
`define ECALL_MI 7'b0101011
`define FENCE_MI 7'b0101100
`define FENCE_I_MI 7'b0101101
`define JAL_MI 7'b0101110
`define JALR_MI 7'b0101111
`define LB_MI 7'b0110000
`define LBU_MI 7'b0110001
`define LH_MI 7'b0110010
`define LHU_MI 7'b0110011
`define LUI_MI 7'b0110100
`define LW_MI 7'b0110101
`define MUL_MI 7'b0110110
`define MULH_MI 7'b0110111
`define MULHSU_MI 7'b0111000
`define MULHU_MI 7'b0111001
`define OR_MI 7'b0111010
`define ORI_MI 7'b0111011
`define REM_MI 7'b0111100
`define REMU_MI 7'b0111101
`define SB_MI 7'b0111110
`define SH_MI 7'b0111111
`define SLL_MI 7'b1000000
`define SLLI_MI 7'b1000001
`define SLT_MI 7'b1000010
`define SLTI_MI 7'b1000011
`define SLTIU_MI 7'b1000100
`define SLTU_MI 7'b1000101
`define SRA_MI 7'b1000110
`define SRAI_MI 7'b1000111
`define SRL_MI 7'b1001000
`define SRLI_MI 7'b1001001
`define SUB_MI 7'b1001010
`define SW_MI 7'b1001011
`define XOR_MI 7'b1001100
`define XORI_MI 7'b1001101

`define HMDST_MI 7'b1001110
`define PKG_MI 7'b1001111
`define RVRS_MI 7'b1010000
`define SLADD_MI 7'b1010001
`define CNTZ_MI 7'b1010010
`define CNTP_MI 7'b1010011

`define CONV_LD_W_MI 7'b1010100
`define CONV_CLR_W_MI 7'b1010101
`define CONV_LD_X_MI 7'b1010110
`define CONV_CLR_X_MI 7'b1010111
`define CONV_RUN_MI 7'b1011000
