
module zero_counter(
    input [31:0] kaynak_yazmac_degeri,
    output reg [4:0] sifir_sayisi,
    output reg [0:0] hepsi_sifir
);
    assign hepsi_sifir = !(|kaynak_yazmac_degeri);
    always@*begin
        case(kaynak_yazmac_degeri)
            32'b00000000_00000000_00000000_00000001:
                sifir_sayisi = 5'd0
            32'b00000000_00000000_00000000_00000010:
                sifir_sayisi = 5'd1
            32'b00000000_00000000_00000000_00000100:
                sifir_sayisi = 5'd2
            32'b00000000_00000000_00000000_00001000:
                sifir_sayisi = 5'd3
            32'b00000000_00000000_00000000_00010000:
                sifir_sayisi = 5'd4
            32'b00000000_00000000_00000000_00100000:
                sifir_sayisi = 5'd5
            32'b00000000_00000000_00000000_01000000:
                sifir_sayisi = 5'd6
            32'b00000000_00000000_00000000_10000000:
                sifir_sayisi = 5'd7
            32'b00000000_00000000_00000001_00000000:
                sifir_sayisi = 5'd8
            32'b00000000_00000000_00000010_00000000:
                sifir_sayisi = 5'd9
            32'b00000000_00000000_00000100_00000000:
                sifir_sayisi = 5'd10
            32'b00000000_00000000_00001000_00000000:
                sifir_sayisi = 5'd11
            32'b00000000_00000000_00010000_00000000:
                sifir_sayisi = 5'd12
            32'b00000000_00000000_00100000_00000000:
                sifir_sayisi = 5'd13
            32'b00000000_00000000_01000000_00000000:
                sifir_sayisi = 5'd14
            32'b00000000_00000000_10000000_00000000:
                sifir_sayisi = 5'd15
            32'b00000000_00000001_00000000_00000000:
                sifir_sayisi = 5'd16
            32'b00000000_00000010_00000000_00000000:
                sifir_sayisi = 5'd17
            32'b00000000_00000100_00000000_00000000:
                sifir_sayisi = 5'd18
            32'b00000000_00001000_00000000_00000000:
                sifir_sayisi = 5'd19
            32'b00000000_00010000_00000000_00000000:
                sifir_sayisi = 5'd20
            32'b00000000_00100000_00000000_00000000:
                sifir_sayisi = 5'd21
            32'b00000000_01000000_00000000_00000000:
                sifir_sayisi = 5'd22
            32'b00000000_10000000_00000000_00000000:
                sifir_sayisi = 5'd23
            32'b00000001_00000000_00000000_00000000:
                sifir_sayisi = 5'd24
            32'b00000010_00000000_00000000_00000000:
                sifir_sayisi = 5'd25
            32'b00000100_00000000_00000000_00000000:
                sifir_sayisi = 5'd26
            32'b00001000_00000000_00000000_00000000:
                sifir_sayisi = 5'd27
            32'b00010000_00000000_00000000_00000000:
                sifir_sayisi = 5'd28
            32'b00100000_00000000_00000000_00000000:
                sifir_sayisi = 5'd29
            32'b01000000_00000000_00000000_00000000:
                sifir_sayisi = 5'd30
            32'b10000000_00000000_00000000_00000000:
                sifir_sayisi = 5'd31
        endcase
    end
endmodule
