// tb_yapay_zeka_hizlandiricisi.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module tb_yapay_zeka_hizlandiricisi();

    yapay_zeka_hizlandiricisi yzh(

    );

    initial begin

        $finish;
    end

endmodule
