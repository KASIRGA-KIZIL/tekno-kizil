// yazmac_obegi.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module yazmac_obegi(
    input clk_i,
    input rst_i


);


endmodule
