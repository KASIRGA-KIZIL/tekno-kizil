// dallanma_ongorucu.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module dallanma_ongorucu(
    input clk_i,
    input rst_i


);


endmodule
