// tb_aritmetik_mantik_birimi.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module tb_aritmetik_mantik_birimi();

    aritmetik_mantik_birimi amb(

    );

    initial begin

        $finish;
    end

endmodule
