// dallanma_birimi.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module dallanma_birimi(


);


endmodule
