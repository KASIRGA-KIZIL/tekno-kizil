// geri_yaz.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module geri_yaz(
    input clk_i,
    input rst_i


);


endmodule
