// pwm_denetleyici.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module pwm_denetleyici(
    input clk_i,
    input rst_i


);


endmodule
