@40000000
B7 07 01 20 13 07 80 09 23 A6 E7 00 37 07 0F 00
13 07 17 00 23 A0 E7 00 37 27 00 00 23 A8 E7 00
37 07 01 20 83 27 47 00 93 F7 27 00 E3 8C 07 FE
93 07 80 09 23 26 F7 00 B7 07 0F 00 93 87 57 00
23 20 F7 00 B7 27 00 00 23 28 F7 00 37 07 01 20
83 27 47 00 93 F7 27 00 E3 8C 07 FE 93 07 80 09
23 26 F7 00 B7 07 0F 00 93 87 97 00 23 20 F7 00
B7 27 00 00 23 28 F7 00 37 07 01 20 83 27 47 00
93 F7 27 00 E3 8C 07 FE 93 07 80 09 23 26 F7 00
B7 07 0F 00 93 87 D7 00 23 20 F7 00 B7 27 00 00
23 28 F7 00 6F 00 00 00
