// modified_booth_dadda_carpici.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module modified_booth_dadda_carpici(


);


endmodule
