// wishbone.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"
// Ornek bus kullanimi icin
module wishbone#(
    parameter SLAVE_SAYISI = 3
)(
    input clk_i,
    input rst_i
    
    
);

endmodule
