@40000000
81 40 01 41 81 41 01 42 81 42 01 43 81 43 01 44
81 44 01 45 81 45 01 46 81 46 01 47 81 47 01 48
81 48 01 49 81 49 01 4A 81 4A 01 4B 81 4B 01 4C
81 4C 01 4D 81 4D 01 4E 81 4E 01 4F 81 4F 85 42
FE 02 63 C8 02 00 05 45 97 12 00 00 23 AC A2 FA
DD BF 97 91 00 00 93 81 61 59 13 82 71 89 13 72
02 FC 13 01 15 00 4A 01 12 91 13 16 25 01 32 92
6F 50 80 25 00 00
@40001000
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00
@40002000
2E 8E 01 48 63 DB 05 00 B3 37 A0 00 33 0E B0 40
33 0E FE 40 33 05 A0 40 7D 58 63 D9 06 00 B3 37
C0 00 B3 06 D0 40 9D 8E 33 06 C0 40 B2 88 AA 87
F2 85 63 9C 06 1A 37 67 00 40 13 07 87 E3 63 7E
CE 0A C1 66 63 74 D6 0A 93 36 06 10 93 C6 16 00
8E 06 33 53 D6 00 1A 97 03 47 07 00 36 97 93 06
00 02 33 83 E6 40 63 8B E6 00 B3 15 6E 00 33 57
E5 00 B3 18 66 00 D9 8D B3 17 65 00 13 D6 08 01
B3 D6 C5 02 13 95 08 01 41 81 13 D7 07 01 B3 F5
C5 02 B3 86 A6 02 C2 05 4D 8F 63 78 D7 00 46 97
63 65 17 01 63 73 D7 00 46 97 15 8F B3 56 C7 02
33 77 C7 02 B3 86 A6 02 C2 07 42 07 C1 83 D9 8F
63 F8 D7 00 C6 97 63 E5 17 01 63 F3 D7 00 C6 97
95 8F 33 D5 67 00 81 45 63 09 08 00 B3 37 A0 00
B3 05 B0 40 9D 8D 33 05 A0 40 82 80 37 03 00 01
C1 46 E3 60 66 F6 E1 46 A9 BF 81 46 09 CA C1 66
63 74 D6 06 93 36 06 10 93 C6 16 00 8E 06 B3 55
D6 00 2E 97 03 47 07 00 36 97 93 06 00 02 33 83
E6 40 63 9A E6 04 33 07 CE 40 93 D5 08 01 33 56
B7 02 13 95 08 01 41 81 93 D6 07 01 33 77 B7 02
33 06 A6 02 42 07 55 8F 63 78 C7 00 46 97 63 65
17 01 63 73 C7 00 46 97 11 8F B3 56 B7 02 33 77
B7 02 B3 86 A6 02 89 BF B7 05 00 01 C1 46 E3 60
B6 FA E1 46 69 BF B3 18 66 00 B3 56 EE 00 B3 17
65 00 33 57 E5 00 13 D5 08 01 B3 D5 A6 02 33 1E
6E 00 33 67 C7 01 13 9E 08 01 13 5E 0E 01 B3 F6
A6 02 B3 85 C5 03 13 96 06 01 93 56 07 01 D1 8E
63 F8 B6 00 C6 96 63 E5 16 01 63 F3 B6 00 C6 96
8D 8E 33 D6 A6 02 42 07 41 83 B3 F6 A6 02 33 06
C6 03 C2 06 55 8F 63 78 C7 00 46 97 63 65 17 01
63 73 C7 00 46 97 11 8F 89 B7 E3 67 DE EE 41 67
63 F6 E6 04 13 B7 06 10 13 47 17 00 0E 07 B7 68
00 40 33 D3 E6 00 93 88 88 E3 9A 98 83 C8 08 00
13 03 00 02 BA 98 33 07 13 41 63 18 13 03 63 E4
C6 01 63 6B C5 00 33 06 C5 40 B3 06 DE 40 B3 35
C5 00 B2 87 B3 85 B6 40 3E 85 79 BD B7 08 00 01
41 47 E3 EE 16 FB 61 47 5D BF B3 96 E6 00 33 53
16 01 33 63 D3 00 B3 57 1E 01 93 5E 03 01 B3 DF
D7 03 33 1E EE 00 B3 55 15 01 B3 E5 C5 01 13 1E
03 01 13 5E 0E 01 33 16 E6 00 33 15 E5 00 B3 F7
D7 03 33 0F FE 03 93 96 07 01 93 D7 05 01 D5 8F
FE 86 63 FC E7 01 9A 97 93 86 FF FF 63 E7 67 00
63 F5 E7 01 93 86 EF FF 9A 97 B3 87 E7 41 33 DF
D7 03 C2 05 C1 81 B3 F7 D7 03 33 0E EE 03 C2 07
DD 8D FA 87 63 FC C5 01 9A 95 93 07 FF FF 63 E7
65 00 63 F5 C5 01 93 07 EF FF 9A 95 C2 06 C1 6F
DD 8E B3 85 C5 41 13 8E FF FF B3 F7 C6 01 93 5E
06 01 C1 82 33 7E C6 01 33 8F C7 03 33 8E C6 03
B3 87 D7 03 B3 86 D6 03 B3 8E C7 01 93 57 0F 01
F6 97 63 F3 C7 01 FE 96 13 DE 07 01 F2 96 41 6E
7D 1E B3 F7 C7 01 C2 07 33 7F CF 01 FA 97 63 E6
D5 00 63 9C D5 00 63 7A F5 00 33 86 C7 40 33 BE
C7 00 B2 87 33 06 6E 00 91 8E B3 07 F5 40 33 35
F5 00 95 8D 89 8D B3 98 15 01 B3 D7 E7 00 33 E5
F8 00 B3 D5 E5 00 8D BB AA 88 2E 83 32 87 2A 88
AE 87 63 96 06 20 B7 65 00 40 93 85 85 E3 63 71
C3 0C C1 66 63 77 D6 0A 93 36 06 10 93 C6 16 00
8E 06 33 55 D6 00 AA 95 83 C5 05 00 13 05 00 02
AE 96 B3 05 D5 40 63 0B D5 00 B3 17 B3 00 B3 D6
D8 00 33 17 B6 00 D5 8F 33 98 B8 00 93 55 07 01
33 D3 B7 02 13 16 07 01 41 82 B3 F7 B7 02 1A 85
B3 08 66 02 93 96 07 01 93 57 08 01 D5 8F 63 FC
17 01 BA 97 13 05 F3 FF 63 E7 E7 00 63 F5 17 01
13 05 E3 FF BA 97 B3 87 17 41 B3 D8 B7 02 42 08
13 58 08 01 B3 F7 B7 02 B3 06 16 03 C2 07 33 68
F8 00 C6 87 63 7B D8 00 3A 98 93 87 F8 FF 63 66
E8 00 63 74 D8 00 93 87 E8 FF 42 05 5D 8D 81 45
82 80 37 05 00 01 C1 46 E3 6D A6 F4 E1 46 91 BF
81 46 09 CA C1 67 63 7F F6 08 93 36 06 10 93 C6
16 00 8E 06 B3 57 D6 00 BE 95 83 C7 05 00 B6 97
93 06 00 02 B3 85 F6 40 63 95 F6 08 B3 07 C3 40
85 45 93 58 07 01 33 DE 17 03 13 16 07 01 41 82
93 56 08 01 B3 F7 17 03 72 85 33 03 C6 03 C2 07
D5 8F 63 FC 67 00 BA 97 13 05 FE FF 63 E7 E7 00
63 F5 67 00 13 05 EE FF BA 97 B3 87 67 40 33 D3
17 03 42 08 13 58 08 01 B3 F7 17 03 B3 06 66 02
C2 07 33 68 F8 00 9A 87 63 7B D8 00 3A 98 93 07
F3 FF 63 66 E8 00 63 74 D8 00 93 07 E3 FF 42 05
5D 8D 82 80 B7 07 00 01 C1 46 E3 65 F6 F6 E1 46
95 B7 33 17 B6 00 B3 56 F3 00 13 55 07 01 33 13
B3 00 B3 D7 F8 00 B3 E7 67 00 33 D3 A6 02 13 16
07 01 41 82 33 98 B8 00 B3 F6 A6 02 B3 08 66 02
93 95 06 01 93 D6 07 01 CD 8E 9A 85 63 FC 16 01
BA 96 93 05 F3 FF 63 E7 E6 00 63 F5 16 01 93 05
E3 FF BA 96 B3 86 16 41 B3 D8 A6 02 C2 07 C1 83
B3 F6 A6 02 33 06 16 03 C2 06 D5 8F C6 86 63 FC
C7 00 BA 97 93 86 F8 FF 63 E7 E7 00 63 F5 C7 00
93 86 E8 FF BA 97 C2 05 91 8F D5 8D DD BD 63 E1
D5 14 C1 67 63 FF F6 02 13 B7 06 10 13 47 17 00
0E 07 B7 67 00 40 B3 D5 E6 00 93 87 87 E3 AE 97
83 C7 07 00 BA 97 13 07 00 02 B3 05 F7 40 63 11
F7 02 05 45 E3 EE 66 E6 33 B5 C8 00 13 45 15 00
82 80 B7 07 00 01 41 47 E3 E5 F6 FC 61 47 D1 B7
33 57 F6 00 B3 96 B6 00 D9 8E 33 57 F3 00 33 13
B3 00 B3 D7 F8 00 B3 E7 67 00 13 D3 06 01 B3 5E
67 02 13 98 06 01 13 58 08 01 33 16 B6 00 33 77
67 02 33 0E D8 03 13 15 07 01 13 D7 07 01 49 8F
76 85 63 7C C7 01 36 97 13 85 FE FF 63 67 D7 00
63 75 C7 01 13 85 EE FF 36 97 33 07 C7 41 33 5E
67 02 C2 07 C1 83 33 77 67 02 33 08 C8 03 42 07
D9 8F 72 87 63 FC 07 01 B6 97 13 07 FE FF 63 E7
D7 00 63 F5 07 01 13 07 EE FF B6 97 42 05 41 6E
59 8D 93 06 FE FF 33 77 D5 00 B3 87 07 41 F1 8E
13 58 05 01 41 82 33 03 D7 02 B3 06 D8 02 33 07
C7 02 33 08 C8 02 33 06 D7 00 13 57 03 01 32 97
63 73 D7 00 72 98 93 56 07 01 C2 96 63 E0 D7 02
E3 97 D7 D8 C1 67 FD 17 7D 8F 42 07 33 73 F3 00
B3 98 B8 00 1A 97 81 45 E3 FC E8 D6 7D 15 85 BB
81 45 01 45 82 80 32 88 AA 87 2E 87 63 93 06 1A
B7 68 00 40 93 88 88 E3 63 F6 C5 0A C1 66 63 7C
D6 08 93 36 06 10 93 C6 16 00 8E 06 33 53 D6 00
9A 98 83 C8 08 00 13 03 00 02 C6 96 B3 08 D3 40
63 0B D3 00 33 97 15 01 B3 56 D5 00 33 18 16 01
55 8F B3 17 15 01 13 56 08 01 B3 56 C7 02 13 15
08 01 41 81 33 77 C7 02 B3 86 A6 02 93 15 07 01
13 D7 07 01 4D 8F 63 78 D7 00 42 97 63 65 07 01
63 73 D7 00 42 97 15 8F B3 56 C7 02 33 77 C7 02
B3 86 A6 02 C2 07 42 07 C1 83 D9 8F 63 F8 D7 00
C2 97 63 E5 07 01 63 F3 D7 00 C2 97 95 8F 33 D5
17 01 81 45 82 80 37 03 00 01 C1 46 E3 68 66 F6
E1 46 AD B7 81 46 09 CA 41 67 63 74 E6 06 93 36
06 10 93 C6 16 00 8E 06 33 57 D6 00 BA 98 03 C7
08 00 36 97 93 06 00 02 B3 88 E6 40 63 9A E6 04
33 87 C5 40 93 55 08 01 33 56 B7 02 13 15 08 01
41 81 93 D6 07 01 33 77 B7 02 33 06 A6 02 42 07
55 8F 63 78 C7 00 42 97 63 65 07 01 63 73 C7 00
42 97 11 8F B3 56 B7 02 33 77 B7 02 B3 86 A6 02
95 B7 37 07 00 01 C1 46 E3 60 E6 FA E1 46 69 BF
33 18 16 01 B3 D6 E5 00 B3 17 15 01 B3 95 15 01
33 57 E5 00 13 55 08 01 4D 8F B3 D5 A6 02 13 13
08 01 13 53 03 01 B3 F6 A6 02 B3 85 65 02 13 96
06 01 93 56 07 01 D1 8E 63 F8 B6 00 C2 96 63 E5
06 01 63 F3 B6 00 C2 96 8D 8E 33 D6 A6 02 42 07
41 83 B3 F6 A6 02 33 06 66 02 C2 06 55 8F 63 78
C7 00 42 97 63 65 07 01 63 73 C7 00 42 97 11 8F
91 B7 63 ED D5 16 41 68 63 F7 06 05 13 B8 06 10
13 48 18 00 0E 08 B7 68 00 40 33 D3 06 01 93 88
88 E3 9A 98 83 C8 08 00 13 03 00 02 C2 98 33 08
13 41 63 19 13 03 63 E4 B6 00 63 6B C5 00 33 06
C5 40 B3 86 D5 40 33 37 C5 00 B2 87 33 87 E6 40
3E 85 BA 85 82 80 B7 08 00 01 41 48 E3 ED 16 FB
61 48 55 BF B3 57 16 01 B3 96 06 01 DD 8E 33 D7
15 01 13 DE 06 01 33 5F C7 03 13 93 06 01 13 53
03 01 B3 97 05 01 B3 55 15 01 DD 8D 93 D7 05 01
33 16 06 01 33 15 05 01 33 77 C7 03 B3 0E E3 03
42 07 D9 8F 7A 87 63 FC D7 01 B6 97 13 07 FF FF
63 E7 D7 00 63 F5 D7 01 13 07 EF FF B6 97 B3 87
D7 41 B3 DE C7 03 C2 05 C1 81 B3 F7 C7 03 76 8E
33 03 D3 03 C2 07 DD 8D 63 FC 65 00 B6 95 13 8E
FE FF 63 E7 D5 00 63 F5 65 00 13 8E EE FF B6 95
93 17 07 01 41 6F B3 E7 C7 01 B3 85 65 40 13 03
FF FF 33 F7 67 00 13 5E 06 01 C1 83 33 73 66 00
B3 0E 67 02 33 83 67 02 33 07 C7 03 B3 87 C7 03
33 0E 67 00 13 D7 0E 01 72 97 63 73 67 00 FA 97
13 53 07 01 9A 97 41 63 7D 13 33 77 67 00 42 07
B3 FE 6E 00 76 97 63 E6 F5 00 63 9B F5 00 63 79
E5 00 33 06 C7 40 33 33 C7 00 9A 96 32 87 95 8F
33 07 E5 40 33 35 E5 00 9D 8D 89 8D B3 98 15 01
33 57 07 01 33 E5 E8 00 B3 D5 05 01 82 80
@400029EE
19 C6 03 15 25 00 83 97 25 00 1D 8D 82 80 83 17
05 00 13 97 07 01 41 83 21 83 93 F7 07 F0 D9 8F
23 10 F5 00 83 97 05 00 03 15 25 00 13 97 07 01
41 83 21 83 93 F7 07 F0 D9 8F 23 90 F5 00 83 97
25 00 1D 8D 82 80
@40002A34
01 11 22 CC 03 14 05 00 06 CE 26 CA 93 57 74 40
4A C8 4E C6 85 8B 91 CB F2 40 13 75 F4 07 62 44
D2 44 42 49 B2 49 05 61 82 80 13 57 34 40 3D 8B
AE 84 93 76 74 00 93 15 47 00 83 D7 84 03 AA 89
D9 8D 95 CE 05 47 63 89 E6 06 13 15 04 01 41 81
22 89 BE 85 EF 10 00 6D AA 87 13 74 04 F0 13 75
F9 07 49 8C 23 9C F4 02 13 64 04 08 23 90 89 00
F2 40 62 44 D2 44 42 49 B2 49 05 61 82 80 93 06
20 02 2E 87 63 D4 D5 00 13 07 20 02 83 96 24 00
03 96 04 00 CC 48 88 4C 13 77 F7 0F EF 10 80 4F
83 D7 E4 03 99 E3 23 9F A4 02 13 19 05 01 83 D7
84 03 13 59 09 41 71 BF 3E 86 13 85 84 02 EF 10
E0 1C 83 D7 C4 03 F5 F3 23 9E A4 02 F9 BF
@40002B02
41 11 26 C2 AE 84 B2 85 06 C6 22 C4 32 84 15 37
AA 87 A2 85 26 85 3E 84 29 3F B2 40 33 05 A4 40
22 44 92 44 41 01 82 80
@40002B2A
03 97 05 00 83 97 25 00 23 10 E5 00 23 11 F5 00
82 80
@40002B3C
03 28 06 00 93 08 88 00 63 FF E8 02 98 42 13 03
47 00 63 7A F3 02 23 20 16 01 1C 41 83 98 05 00
03 96 25 00 23 20 F8 00 23 20 05 01 23 22 E8 00
9C 42 42 85 91 07 9C C2 83 27 48 00 23 90 17 01
23 91 C7 00 82 80 01 48 42 85 82 80
@40002B88
AA 87 08 41 D4 43 50 41 18 41 D0 C3 54 C1 98 C3
23 20 05 00 82 80
@40002B9E
D0 41 54 41 98 41 50 C1 D4 C1 18 C1 88 C1 82 80
@40002BAE
03 97 25 00 63 4C 07 00 01 E5 3D A0 08 41 1D C1
5C 41 83 97 27 00 E3 9B E7 FE 82 80 01 CD 03 97
05 00 19 A0 08 41 01 C9 5C 41 83 C7 07 00 E3 9B
E7 FE 82 80 01 45 82 80 82 80
@40002BE8
01 C9 01 47 11 A0 3E 85 1C 41 18 C1 2A 87 E5 FF
82 80
@40002BFA
79 71 4E CE 56 CA 5E C6 62 C4 6A C0 06 D6 22 D4
26 D2 4A D0 52 CC 5A C8 66 C2 AA 89 2E 8C B2 8B
85 4A 05 4D 63 83 09 08 81 4C 81 44 01 4B 85 0C
CE 87 01 44 9C 43 05 04 99 C3 E3 9D 8A FE 4E 89
56 8A BE 89 63 5D 80 00 63 18 0A 02 CA 87 03 29
09 00 7D 14 99 CC 9C C0 BE 84 E3 47 80 FE 63 5C
40 03 63 8C 09 02 19 E8 CE 87 7D 1A 83 A9 09 00
FD F0 3E 8B BE 84 D5 B7 E3 8A 09 FC 83 A5 49 00
03 25 49 00 5E 86 02 9C E3 52 A0 FC CE 87 7D 1A
83 A9 09 00 C1 B7 E3 9C 09 F8 23 A0 04 00 63 89
AC 01 DA 89 86 0A E3 91 09 F8 23 20 00 00 02 90
B2 50 22 54 92 54 02 59 F2 49 62 4A D2 4A B2 4B
22 4C 92 4C 02 4D 5A 85 42 4B 45 61 82 80
@40002CC8
2A 86 03 15 45 00 01 11 22 CC 26 CA 06 CE 4A C8
4E C6 52 C4 56 C2 40 52 AE 84 63 5D A0 1A 81 48
01 4E 01 43 01 48 13 FA F8 0F 63 CA 04 14 63 06
04 1A A2 87 19 A0 9C 43 91 C7 D8 43 03 17 27 00
E3 1B 97 FE 81 46 11 A0 3A 84 18 40 14 C0 A2 86
65 FF 63 82 07 14 D8 43 03 17 07 00 93 76 17 00
81 CA 25 87 05 8B 42 97 13 18 07 01 13 58 08 01
98 43 11 C7 14 43 94 C3 1C 40 1C C3 18 C0 05 03
42 03 13 53 03 01 63 C5 04 00 85 04 C2 04 C1 84
85 08 C2 08 93 D8 08 41 E3 17 15 F9 93 17 23 00
B3 87 C7 41 3E 98 13 19 08 01 13 59 09 01 63 59
B0 00 22 85 97 05 00 00 93 85 65 D8 9D 3D 2A 84
1C 40 A2 89 83 AA 07 00 D8 43 03 A6 4A 00 83 A6
0A 00 D0 C3 23 A2 EA 00 94 C3 23 A0 0A 00 63 D7
04 00 79 A0 83 A9 09 00 63 86 09 0C 83 A7 49 00
83 97 27 00 E3 98 97 FE 5C 40 CA 85 03 95 07 00
EF 10 20 49 83 A9 09 00 2A 89 E3 97 09 FE 83 29
04 00 03 A7 4A 00 83 A6 49 00 83 A7 09 00 22 85
23 A2 DA 00 23 A2 E9 00 23 A0 FA 00 01 46 23 A0
59 01 97 05 00 00 93 85 45 BF E5 3B 00 41 AA 84
11 C8 DC 40 CA 85 03 95 07 00 EF 10 80 44 00 40
2A 89 65 F8 F2 40 62 44 D2 44 B2 49 22 4A 92 4A
4A 85 42 49 05 61 82 80 83 A9 09 00 63 84 09 04
83 A7 49 00 83 C7 07 00 E3 18 FA FE B5 BF 31 CC
A2 87 21 A0 9C 43 E3 8F 07 EA D8 43 03 47 07 00
E3 1A EA FE 45 BD 1C 40 05 0E 42 0E DC 43 13 5E
0E 01 83 87 17 00 85 8B C2 97 13 98 07 01 13 58
08 01 D1 BD 83 29 04 00 E3 8F 09 F4 5C 40 CA 85
03 95 07 00 EF 10 E0 3C 83 A9 09 00 2A 89 E3 95
09 F2 35 BF 01 49 01 4A D9 BD 83 27 00 00 02 90
@40002EA8
D1 47 33 5E F5 02 E1 77 23 A0 05 00 13 87 07 08
93 86 05 01 2E 85 13 83 85 00 79 1E 13 1F 3E 00
2E 9F 23 A2 E5 01 93 1F 2E 00 23 10 EF 00 23 11
0F 00 FA 9F 13 07 4F 00 63 FC E6 0F 93 08 8F 00
63 F8 F8 0F D8 C5 23 A4 05 00 23 A0 65 00 93 C7
F7 FF 7D 57 23 12 EF 00 23 13 FF 00 63 0E 0E 04
93 12 06 01 E1 73 93 D2 02 01 01 48 93 C3 F3 FF
13 17 08 01 41 83 B3 C7 E2 00 8E 07 1D 8B 93 F7
87 07 D9 8F 13 97 87 00 93 85 86 00 05 08 93 8E
48 00 5D 8F 63 F0 E5 03 63 FE FE 01 23 A0 66 00
14 C1 23 A2 16 01 23 90 E8 00 23 91 78 00 36 83
F6 88 AE 86 E3 1E 0E FB 03 28 03 00 63 04 08 06
95 47 91 6E 33 5E FE 02 13 07 00 20 85 46 FD 1E
0D A0 93 97 06 01 83 28 08 00 C1 87 13 07 07 10
42 07 23 91 F5 00 42 83 85 06 41 83 63 8C 08 02
46 88 B3 C5 C6 00 93 77 07 70 CD 8F B3 F7 D7 01
83 25 43 00 E3 E7 C6 FD 83 28 08 00 C2 07 C1 87
13 07 07 10 42 07 23 91 F5 00 42 83 85 06 41 83
E3 98 08 FC 01 46 97 05 00 00 93 85 05 A2 15 B1
9A 86 BA 88 01 43 1D B7
@40002FE0
41 11 4A C0 03 29 C5 01 06 C6 22 C4 26 C2 23 2C
05 02 23 2E 05 02 63 0C 09 02 2A 84 81 44 85 45
22 85 D9 31 83 55 84 03 EF 10 00 15 FD 55 23 1C
A4 02 22 85 55 39 83 55 84 03 EF 10 E0 13 23 1C
A4 02 99 E0 23 1D A4 02 85 04 E3 1A 99 FC B2 40
22 44 92 44 02 49 01 45 41 01 82 80
@4000303C
FD 77 05 67 19 71 93 87 C7 7D 13 07 07 83 86 DE
3E 97 A2 DC A6 DA CA D8 CE D6 D2 D4 D6 D2 DA D0
DE CE E2 CC E6 CA EA C8 EE C6 13 01 01 81 2E 86
2A C6 B3 05 27 00 13 05 E1 05 EF 10 60 2D 17 25
00 00 13 05 65 3E EF 10 A0 4D 05 45 EF 10 C0 05
AA 87 09 45 23 1E F1 00 EF 10 00 05 AA 87 0D 45
23 1F F1 00 EF 10 40 04 AA 87 11 45 23 10 F1 02
EF 10 80 03 AA 87 15 45 3E DC EF 10 E0 02 11 E1
1D 45 05 67 FD 77 13 07 07 83 3E 97 B3 07 27 00
3E C4 83 A7 C7 7E 2A DE 63 91 07 56 A2 47 83 97
07 7F 63 87 07 58 85 65 FD 76 93 85 05 83 B6 95
B3 86 25 00 90 10 93 77 25 00 13 77 15 00 B3 37
F0 00 36 C4 23 AA C6 7E 23 1E 01 04 93 76 45 00
3E 97 81 C6 05 07 42 07 41 83 93 06 00 7D B3 D6
E6 02 FD 77 05 67 93 87 C7 7E 13 07 07 83 3E 97
B3 07 27 00 01 48 01 47 05 43 8D 48 36 DA B3 15
E3 00 E9 8D 05 07 63 91 05 4E 91 07 E3 19 17 FF
85 66 7D 77 F2 57 93 86 06 83 BA 96 33 87 26 00
3A C4 13 F7 17 00 11 CB A2 47 52 55 03 96 C7 7E
83 A5 87 7F 25 3B F2 57 AA C0 13 F7 27 00 63 11
07 20 91 8B 99 CF 05 67 FD 77 13 07 07 83 3E 97
B3 07 27 00 42 56 83 95 C7 7E 52 55 3E C4 EF 00
50 34 E2 57 A9 E7 85 47 7D 74 3E DC 85 67 13 04
C4 7E 93 87 07 83 A2 97 33 84 27 00 62 57 93 17
27 00 BA 97 86 07 3E DC EF 10 80 12 22 85 19 3D
EF 10 60 13 EF 10 80 14 EF 10 A0 16 65 D1 A9 47
B3 D7 A7 02 62 57 85 07 B3 87 E7 02 3E DC EF 10
20 10 7D 74 85 64 13 05 C4 7E 93 87 04 83 AA 97
33 85 27 00 C5 33 EF 10 00 10 EF 10 20 11 93 87
04 83 A2 97 8A 97 AA 89 03 95 C7 7E 2E 8A 81 45
3E C4 EF 10 C0 03 A2 47 AA 85 03 95 E7 7E EF 10
00 03 A2 47 AA 85 03 95 07 7F EF 10 40 02 AA 85
03 15 41 03 EF 10 A0 01 A1 67 93 87 57 B0 2A 89
63 0C F5 46 63 EB A7 16 89 67 93 87 27 8F 63 05
F5 48 95 67 93 87 F7 EA 63 18 F5 48 17 25 00 00
13 05 05 26 EF 10 C0 2E 89 47 17 6C 00 00 13 0C
2C B7 03 27 0C 00 63 04 07 16 05 67 FD 76 13 07
07 83 36 97 86 07 0A 97 97 2D 00 00 93 8D CD 7C
81 4A 81 4C 3A C4 05 6D BE 9D 97 2B 00 00 93 8B
2B 2B 17 2B 00 00 13 0B AB 2D 0D A8 22 47 B3 07
94 01 8A 07 BA 97 EA 97 83 D7 C7 82 85 0C 83 26
0C 00 D6 97 C2 0C 93 94 07 01 93 9A 07 01 93 DC
0C 01 C1 80 93 DA 0A 41 63 F4 DC 10 A2 47 13 94
4C 00 B3 04 94 01 8A 04 BE 94 EA 94 83 A7 C4 80
23 96 04 82 93 F6 17 00 95 C2 03 D6 64 82 83 D6
0D 00 63 0D D6 00 E6 85 5E 85 EF 10 60 24 83 D6
C4 82 83 A7 C4 80 85 06 23 96 D4 82 93 F6 27 00
85 CA 22 47 B3 04 94 01 8A 04 BA 94 EA 94 03 D6
84 82 83 D6 CD 00 63 0D D6 00 E6 85 5A 85 EF 10
20 21 83 D6 C4 82 83 A7 C4 80 85 06 23 96 D4 82
91 8B A9 DF A2 47 66 94 0A 04 3E 94 6A 94 03 56
A4 82 83 D6 8D 01 63 1B D6 02 83 57 C4 82 B9 B7
05 67 FD 77 13 07 07 83 3E 97 B3 07 27 00 3E C4
22 47 83 97 E7 7E 52 55 03 16 C7 7E 83 25 C7 7F
C2 07 5D 8E D4 00 AD 2E F2 57 E1 BB E6 85 17 25
00 00 13 05 25 21 EF 10 A0 1A 83 57 C4 82 85 07
C2 07 C1 83 23 16 F4 82 11 B7 A5 67 93 87 27 A0
63 04 F5 30 BD 67 93 87 57 9F 63 1F F5 30 17 25
00 00 13 05 25 12 EF 10 A0 17 8D 47 79 B5 81 44
EF 00 B0 6C D2 55 AA 94 17 25 00 00 13 05 85 1F
EF 10 00 16 CE 85 17 25 00 00 13 05 25 20 EF 10
20 15 D2 85 4E 85 EF 00 D0 72 AA 85 17 25 00 00
13 05 45 20 EF 10 C0 13 C2 04 4E 85 D2 85 C1 80
EF 00 30 71 63 13 05 26 4E 85 D2 85 EF 00 70 70
A5 47 63 F4 A7 24 83 27 0C 00 E2 55 17 25 00 00
13 05 45 24 C2 04 B3 85 F5 02 C1 84 EF 10 40 10
97 25 00 00 93 85 85 24 17 25 00 00 13 05 C5 24
EF 10 00 0F 97 25 00 00 93 85 85 25 17 25 00 00
13 05 05 30 EF 10 C0 0D 97 25 00 00 93 85 C5 30
17 25 00 00 13 05 C5 30 EF 10 80 0C CA 85 17 25
00 00 13 05 65 31 EF 10 A0 0B F2 57 13 F7 17 00
39 C7 03 27 0C 00 21 C7 05 67 FD 77 13 07 07 83
3E 97 B3 07 27 00 01 44 3E C4 85 69 17 29 00 00
13 09 49 30 22 47 93 17 44 00 A2 97 8A 07 BA 97
CE 97 03 D6 67 82 A2 85 4A 85 EF 10 60 07 05 04
83 27 0C 00 42 04 41 80 E3 6E F4 FC F2 57 13 F7
27 00 21 CB 03 27 0C 00 63 0C 07 1A 05 67 FD 77
13 07 07 83 3E 97 B3 07 27 00 01 44 3E C4 85 69
17 29 00 00 13 09 C9 2C 22 47 93 17 44 00 A2 97
8A 07 BA 97 CE 97 03 D6 87 82 A2 85 4A 85 EF 10
20 02 05 04 83 27 0C 00 42 04 41 80 E3 6E F4 FC
F2 57 91 8B 03 27 0C 00 A1 C7 01 44 59 C7 05 67
FD 77 13 07 07 83 3E 97 B3 07 27 00 3E C4 85 69
17 29 00 00 13 09 89 29 22 47 93 17 44 00 A2 97
8A 07 BA 97 CE 97 03 D6 A7 82 A2 85 4A 85 EF 00
30 7D 05 04 83 27 0C 00 42 04 41 80 E3 6E F4 FC
83 27 0C 00 01 44 B1 C3 05 67 FD 77 13 07 07 83
3E 97 B3 07 27 00 3E C4 85 69 17 29 00 00 13 09
A9 26 22 47 93 17 44 00 A2 97 8A 07 BA 97 CE 97
03 D6 47 82 A2 85 4A 85 EF 00 90 78 05 04 83 27
0C 00 42 04 41 80 E3 6E F4 FC C9 C8 63 4B 90 06
17 25 00 00 13 05 C5 29 EF 00 90 76 13 05 E1 05
EF 00 50 56 13 01 01 7F F6 50 66 54 D6 54 46 59
B6 59 26 5A 96 5A 06 5B F6 4B 66 4C D6 4C 46 4D
B6 4D 01 45 09 61 82 80 B3 05 D8 02 05 08 42 08
13 58 08 01 B2 95 CC C7 09 BE 05 47 E3 95 E7 AA
A2 47 83 97 07 7F E3 90 07 AA 22 47 B7 37 15 34
93 87 57 41 23 26 F7 7E 93 07 60 06 23 18 F7 7E
59 B4 17 25 00 00 13 05 E5 28 EF 00 70 6F 79 B7
22 47 93 07 60 06 23 18 F7 7E B5 B4 17 25 00 00
13 05 45 1C EF 00 D0 6D 95 BF 17 25 00 00 13 05
65 FC EF 00 F0 6C 85 04 7D B3 83 27 0C 00 62 54
D2 85 4E 85 33 04 F4 02 EF 00 B0 49 AA 85 17 25
00 00 13 05 A5 F8 B3 55 B4 02 EF 00 70 6A AD BB
91 8B E3 8F 07 EC 15 B7 17 25 00 00 13 05 85 DD
EF 00 10 69 85 47 55 B6 17 25 00 00 13 05 85 D9
EF 00 10 68 81 47 51 BE 17 25 00 00 13 05 85 E4
EF 00 10 67 91 47 51 B6 41 64 93 04 F4 FF 17 5C
00 00 13 0C EC 6E ED B1 41 11 17 25 00 00 13 05
65 33 06 C6 EF 10 F0 1E B2 40 7D 55 41 01 82 80
@4000371C
41 11 22 C6 26 C4 4A C2 4E C0 2A 88 11 E2 05 46
81 47 63 08 08 0A 3E 85 85 07 33 87 F7 02 0E 07
E3 6B 07 FF B3 02 A5 02 FD 15 93 F7 C5 FF 93 84
47 00 2A 89 26 8E 86 02 B3 83 54 00 35 C1 C1 6E
13 03 15 00 13 14 15 00 1E 8F 81 4F 05 47 33 0E
7E 40 FD 1E BA 89 7A 88 33 06 E6 02 93 17 07 01
C1 83 B3 08 0E 01 09 08 05 07 93 55 F6 41 C1 81
2E 96 33 76 D6 01 0D 8E B3 85 C7 00 C2 05 C1 81
AE 97 23 1F B8 FE 93 F7 F7 0F 23 90 F8 00 E3 15
67 FC 85 0F 33 07 35 01 2A 93 22 9F E3 9C AF FA
B3 87 53 00 FD 17 32 44 F1 9B 91 07 C4 C2 23 A0
26 01 23 A4 76 00 DC C6 A2 44 12 49 82 49 41 01
82 80 FD 15 93 F3 C5 FF 13 8E 43 00 F2 84 99 03
7D 59 89 42 7D 55 A5 B7
@400037F4
AA 8E 31 CD 93 1F 25 00 33 0F A0 40 B3 88 F5 01
01 4E 01 45 01 47 81 45 0E 0F 33 83 F8 41 9A 87
31 A0 42 05 91 07 41 85 63 85 F8 02 BA 86 98 43
42 05 41 81 B3 A6 E6 00 BA 95 13 08 A5 00 36 95
E3 51 B6 FE 13 15 08 01 91 07 41 85 81 45 E3 9F
F8 FC 05 0E B3 08 E3 41 E3 91 CE FD 82 80 01 45
82 80
@40003856
21 C1 13 1F 15 00 B3 0E A0 40 33 08 E6 01 01 43
01 4E 8A 0E B3 08 E8 41 13 16 23 00 2E 96 C6 87
03 97 07 00 11 06 89 07 33 07 D7 02 23 2E E6 FE
E3 18 F8 FE 05 0E 2A 93 33 88 D8 41 E3 1C C5 FD
82 80
@40003898
1D C9 13 13 15 00 B3 08 A0 40 42 06 41 82 B3 86
65 00 01 48 8A 08 B3 85 66 40 AE 87 03 D7 07 00
89 07 32 97 23 9F E7 FE E3 9A F6 FE 05 08 B3 86
15 41 E3 12 05 FF 82 80
@400038D0
15 CD 13 1F 25 00 13 1E 15 00 2E 9F 36 9E 81 4E
13 98 1E 00 32 98 B6 87 81 48 03 17 08 00 03 93
07 00 89 07 09 08 33 07 67 02 BA 98 E3 17 FE FE
23 A0 15 01 91 05 AA 9E E3 1C BF FC 82 80
@4000390E
2D C5 41 11 2A 8F 06 05 22 C6 AE 83 36 84 B2 8E
33 08 A6 00 81 4F 81 42 93 98 2F 00 9E 98 22 83
01 4E 9A 86 F6 87 01 46 03 97 07 00 83 95 06 00
89 07 AA 96 33 07 B7 02 3A 96 E3 17 F8 FE 23 A0
C8 00 93 07 1E 00 91 08 09 03 63 04 FF 00 3E 8E
C9 BF 93 87 12 00 AA 9E FA 9F 2A 98 63 84 C2 01
BE 82 5D BF 32 44 41 01 82 80 82 80
@4000397A
2D CD 41 11 2A 8F 06 05 22 C6 AE 83 36 84 B2 8E
33 08 A6 00 81 4F 81 42 93 98 2F 00 9E 98 22 83
01 4E 1A 86 F6 86 81 45 03 17 06 00 83 97 06 00
89 06 2A 96 B3 87 E7 02 13 D7 27 40 95 87 3D 8B
93 F7 F7 07 B3 07 F7 02 BE 95 E3 1F D8 FC 23 A0
B8 00 93 07 1E 00 91 08 09 03 63 04 FF 00 3E 8E
C9 B7 93 87 12 00 AA 9E FA 9F 2A 98 63 84 C2 01
BE 82 5D B7 32 44 41 01 82 80 82 80
@400039F6
39 71 22 DC 26 DA 5A D0 06 DE 4A D8 4E D6 52 D4
56 D2 5E CE 62 CC 66 CA 6A C8 6E C6 2E 8B 32 84
B6 84 63 05 05 24 13 1F 15 00 B3 05 E6 01 B3 0C
A0 40 93 19 07 01 AA 8D 93 D9 09 01 2E 86 01 48
93 98 2C 00 33 03 E6 41 9A 87 83 D6 07 00 89 07
CE 96 23 9F D7 FE E3 9A C7 FE 13 05 18 00 33 06
13 41 63 84 AD 00 2A 88 F1 BF 01 4E 81 4E 33 83
E5 41 13 16 2E 00 5A 96 9A 87 83 96 07 00 11 06
89 07 B3 86 E6 02 23 2E D6 FE E3 98 F5 FE 93 87
1E 00 2A 9E B3 05 13 41 63 84 0E 01 BE 8E C1 BF
33 0E A0 40 FD 77 33 69 F7 00 33 03 1B 41 01 45
01 47 01 46 01 4F 0E 0E B3 0E 13 01 F6 87 31 A0
42 05 91 07 41 85 63 85 67 02 BA 86 98 43 42 05
41 81 B3 A6 E6 00 3A 96 93 05 A5 00 36 95 E3 51
C9 FE 13 95 05 01 91 07 41 85 01 46 E3 9F 67 FC
93 07 1F 00 33 83 CE 41 63 04 E8 01 3E 8F 6D BF
81 45 EF 00 20 76 22 86 AA 8B A6 86 6E 85 DA 85
13 9A 2D 00 D9 33 5A 9A 13 9C 2C 00 52 88 01 45
01 47 01 46 81 4A 8E 0C B3 08 0C 01 C6 87 31 A0
42 05 91 07 41 85 63 85 07 03 BA 86 98 43 42 05
41 81 B3 A6 E6 00 3A 96 93 05 A5 00 36 95 E3 51
C9 FE 13 95 05 01 91 07 41 85 01 46 E3 9F 07 FD
13 8D 1A 00 33 88 98 41 63 84 AD 01 EA 8A 6D BF
DE 85 EF 00 20 6F 22 86 AA 8B A6 86 6A 85 DA 85
61 3B 52 88 01 45 01 47 01 46 01 43 B3 08 88 01
C6 87 31 A0 42 05 91 07 41 85 63 05 F8 02 BA 86
98 43 42 05 41 81 B3 A6 E6 00 3A 96 93 05 A5 00
36 95 E3 51 C9 FE 13 95 05 01 91 07 41 85 01 46
E3 1F F8 FC 93 07 13 00 33 88 98 41 63 04 53 01
3E 83 6D BF DE 85 EF 00 E0 68 AA 87 A6 86 22 86
6A 85 DA 85 BE 84 79 3B 01 45 01 47 01 46 81 48
33 08 8A 01 C2 87 31 A0 42 05 91 07 41 85 63 05
FA 02 BA 86 98 43 42 05 41 81 B3 A6 E6 00 3A 96
93 05 A5 00 36 95 E3 51 C9 FE 13 95 05 01 91 07
41 85 01 46 E3 1F FA FC 93 87 18 00 33 0A 98 41
63 84 58 01 BE 88 6D BF A6 85 EF 00 A0 62 06 0D
6A 94 01 46 B3 06 A4 41 B6 87 03 D7 07 00 89 07
33 07 37 41 23 9F E7 FE E3 99 87 FE 93 07 16 00
33 84 86 41 63 02 56 05 3E 86 E9 BF 81 45 DD 2B
22 86 2A 89 A6 86 01 45 DA 85 85 31 CA 85 01 45
D5 23 22 86 A6 86 2A 89 DA 85 01 45 71 31 CA 85
01 45 C9 2B AA 87 22 86 01 45 DA 85 A6 86 3E 84
D5 31 A2 85 01 45 7D 2B F2 50 62 54 42 05 D2 54
42 59 B2 59 22 5A 92 5A 02 5B F2 4B 62 4C D2 4C
42 4D B2 4D 41 85 21 61 82 80
@40003CC0
41 11 22 C4 14 45 32 84 2E 87 50 41 4C 45 08 41
06 C6 15 33 A2 85 22 44 B2 40 41 01 BD AB
@40003CDE
13 08 F5 FF 85 47 63 F2 07 0D 85 05 C2 05 C1 81
41 11 93 D7 35 00 22 C6 1D 4E 93 F6 75 00 01 47
97 2E 00 00 93 8E 6E D8 11 43 85 48 13 0F C0 02
8D 8B 63 8D C6 05 63 65 D3 08 F5 16 C2 06 8A 07
C1 82 F6 97 63 EB D8 06 9C 4B A1 42 93 06 17 00
33 84 56 00 63 76 04 05 32 97 BA 86 B3 83 57 00
83 CF 07 00 85 07 85 06 A3 8F F6 FF E3 9A F3 FE
85 05 C2 05 16 97 C1 81 23 00 E7 01 93 D7 35 00
93 F6 75 00 22 87 8D 8B E3 97 C6 FB 8A 07 A1 42
93 06 17 00 F6 97 33 84 56 00 9C 5B E3 6E 04 FB
63 64 A7 00 01 A8 85 06 32 97 23 00 07 00 36 87
E3 EB A6 FE 32 44 41 01 82 80 9C 43 91 42 79 B7
8A 07 F6 97 9C 53 A1 42 51 B7 01 47 85 46 11 A0
85 06 32 97 23 00 07 00 36 87 E3 EB A6 FE 82 80
@40003DBE
18 41 2A 86 83 46 07 00 63 85 06 1C 93 07 C0 02
01 45 63 80 F6 16 13 85 06 FD 13 75 F5 0F 25 48
63 78 A8 02 13 05 D0 02 63 8E A6 14 13 05 E0 02
63 86 A6 06 13 05 B0 02 63 86 A6 14 D4 41 9C 41
05 07 85 06 85 07 D4 C1 9C C1 05 45 18 C2 82 80
88 41 93 06 17 00 05 05 88 C1 03 47 17 00 63 04
07 16 63 06 F7 10 93 07 E0 02 63 0E F7 0E 13 07
07 FD 13 77 F7 0F A5 47 63 EA E7 00 03 C7 16 00
85 06 63 02 07 14 93 07 C0 02 E1 BF 9C 49 13 87
16 00 05 45 85 07 9C C9 18 C2 82 80 88 41 93 06
17 00 05 05 88 C1 03 47 17 00 63 01 07 12 63 03
F7 14 93 77 F7 0D 13 05 50 04 63 80 A7 02 13 07
07 FD 13 77 F7 0F A5 47 63 E7 E7 0A 03 C7 16 00
85 06 6D CF 93 07 C0 02 D9 BF DC 49 13 87 16 00
85 07 DC C9 83 C7 16 00 ED CB 13 05 C0 02 63 88
A7 0E D8 45 93 87 57 FD 93 F7 D7 0F 05 07 D8 C5
91 C7 13 87 26 00 05 45 18 C2 82 80 83 C7 26 00
13 87 26 00 E9 C3 63 87 A7 0C 88 4D 93 87 07 FD
93 F7 F7 0F 05 05 25 48 88 CD 63 77 F8 00 13 87
36 00 05 45 18 C2 82 80 25 45 83 46 17 00 3A 88
93 08 C0 02 93 87 06 FD 05 07 93 F7 F7 0F CD C2
63 8D 16 09 E3 73 F5 FE DC 41 13 07 28 00 05 45
85 07 DC C1 15 BF 9C 49 85 07 9C C9 85 B7 36 87
11 45 05 07 15 B7 DC 49 13 87 16 00 05 45 85 07
DC C9 19 BF 88 41 93 06 17 00 05 05 88 C1 03 48
17 00 63 09 08 06 63 03 F8 06 98 45 93 07 08 FD
93 F7 F7 0F 25 45 05 07 63 7B F5 00 93 07 E0 02
63 09 F8 00 98 C5 05 45 13 87 16 00 F1 BD 98 C5
75 BD 98 C5 21 B7 36 87 11 45 F9 B5 36 87 15 45
E1 B5 01 45 D1 B5 19 45 C1 B5 0D 45 75 BD 0D 45
05 07 5D BD 19 45 05 07 45 BD 1D 45 05 07 6D B5
1D 45 5D B5 36 87 15 45 05 07 79 BD 36 87 09 45
05 07 59 BD 36 87 09 45 41 BD
@40003FC8
19 71 A6 DA CE D6 04 08 93 09 01 03 A2 DC CA D8
D2 D4 DA D0 DE CE E2 CC 36 8B 3A 8A 3E 89 86 DE
D6 D2 2E 84 2A 8C B2 8B 2E C6 94 08 26 87 CE 87
23 A0 07 00 23 20 07 00 91 07 11 07 E3 9A D7 FE
83 47 04 00 93 0A C1 00 F1 C7 0C 18 56 85 65 33
13 18 25 00 93 07 08 05 33 88 27 00 32 47 83 27
08 FC 03 47 07 00 85 07 23 20 F8 FC 79 FF 22 C6
22 9C 63 75 84 03 A2 87 13 06 C0 02 03 C7 07 00
B3 46 77 01 63 04 C7 00 23 80 D7 00 D2 97 E3 E7
87 FF 83 47 04 00 93 0A C1 00 9D C3 0C 18 56 85
99 3B 13 16 25 00 93 07 06 05 33 86 27 00 32 47
83 27 06 FC 03 47 07 00 85 07 23 20 F6 FC 79 FF
22 C6 93 06 C0 02 63 7D 84 01 83 47 04 00 33 C7
67 01 63 84 D7 00 23 00 E4 00 52 94 E3 67 84 FF
13 84 04 02 88 40 CA 85 91 04 ED 28 AA 85 03 A5
09 00 91 09 C5 28 2A 89 E3 16 94 FE F6 50 66 54
D6 54 46 59 B6 59 26 5A 96 5A 06 5B F6 4B 66 4C
09 61 82 80 22 9C E3 60 84 F7 D9 B7
@400040E4
95 47 63 E2 A7 04 17 27 00 00 13 07 A7 9D 0A 05
3A 95 1C 41 BA 97 82 87 17 55 00 00 03 25 C5 D0
82 80 17 55 00 00 03 25 A5 D0 82 80 17 55 00 00
03 25 C5 CF 82 80 03 A5 81 80 82 80 17 55 00 00
03 25 C5 CC 82 80 01 45 82 80
@4000412E
AA 86 2E 85 E9 75 A1 47 85 05 33 C7 A6 00 FD 17
05 81 05 8B 93 F7 F7 0F 33 46 B5 00 85 82 01 C7
13 15 06 01 41 81 F5 F3 82 80
@40004158
AA 86 69 78 2E 85 13 F6 F6 0F A1 47 05 08 33 47
A6 00 FD 17 05 81 05 8B 93 F7 F7 0F B3 45 05 01
05 82 01 C7 13 95 05 01 41 81 F5 F3 E9 75 A1 82
A1 47 85 05 33 C7 A6 00 FD 17 05 81 05 8B 93 F7
F7 0F 33 46 B5 00 85 82 01 C7 13 15 06 01 41 81
F5 F3 82 80
@400041AC
2A 87 13 16 07 01 E9 78 2E 85 41 82 93 75 F7 0F
A1 47 85 08 B3 C6 A5 00 FD 17 05 81 85 8A 93 F7
F7 0F 33 48 15 01 85 81 81 C6 13 15 08 01 41 81
F5 F3 69 78 21 82 A1 47 05 08 B3 46 A6 00 FD 17
05 81 85 8A 93 F7 F7 0F B3 45 05 01 05 82 81 C6
13 95 05 01 41 81 F5 F3 13 56 07 01 69 78 32 87
A1 47 13 76 F6 0F 05 08 B3 46 A6 00 FD 17 05 81
85 8A 93 F7 F7 0F B3 45 05 01 05 82 81 C6 13 95
05 01 41 81 F5 F3 E9 75 21 83 A1 47 85 05 B3 46
A7 00 FD 17 05 81 85 8A 93 F7 F7 0F 33 46 B5 00
05 83 81 C6 13 15 06 01 41 81 F5 F3 82 80
@4000425A
AA 86 13 96 06 01 69 78 2E 85 41 82 93 F6 F6 0F
A1 47 05 08 33 C7 A6 00 FD 17 05 81 05 8B 93 F7
F7 0F B3 45 05 01 85 82 01 C7 13 95 05 01 41 81
F5 F3 E9 75 93 56 86 00 A1 47 85 05 33 C7 A6 00
FD 17 05 81 05 8B 93 F7 F7 0F 33 46 B5 00 85 82
01 C7 13 15 06 01 41 81 F5 F3 82 80
@400042B6
01 45 82 80
@400042BA
B7 07 08 02 85 07 37 07 00 20 1C C3 82 80
@400042C8
B7 07 00 30 88 43 82 80
@400042D0
B7 07 00 30 C8 43 81 45 82 80
@400042DA
B7 07 00 30 88 43 82 80
@400042E2
B7 07 00 30 CC 43 88 43 82 80
@400042EC
B7 07 00 30 D4 43 98 43 97 57 00 00 93 87 C7 B0
D4 C3 98 C3 82 80
@40004302
B7 07 00 30 D4 43 98 43 97 57 00 00 93 87 E7 AE
D4 C3 98 C3 82 80
@40004318
97 56 00 00 93 86 06 AE 17 57 00 00 13 07 07 AE
9C 42 08 43 CC 42 58 43 33 85 A7 40 B3 B7 A7 00
99 8D 9D 8D 82 80
@4000433E
B7 87 93 03 93 87 07 70 33 55 F5 02 82 80
@4000434C
B7 07 08 02 85 07 37 07 00 20 1C C3 85 47 23 00
F5 00 82 80
@40004360
23 00 05 00 82 80
@40004366
1D 71 A2 CE A6 CC 13 F8 07 04 97 1E 00 00 93 8E
0E 68 63 16 08 00 97 1E 00 00 93 8E CE 64 13 F4
07 01 63 14 04 10 13 F8 17 00 93 F4 17 01 93 03
00 03 63 0E 08 0E 13 F8 27 00 13 FF 07 02 63 04
08 0E 63 CF 05 0E 13 F8 47 00 63 17 08 12 A1 8B
81 4F 81 C7 FD 16 93 0F 00 02 63 0A 0F 00 C1 47
63 00 F6 14 93 07 86 FF 93 B7 17 00 9D 8E E5 E1
93 07 00 03 23 06 F1 00 05 48 93 02 C1 00 C2 88
63 53 E8 00 BA 88 B3 86 16 41 89 EC 33 07 D5 00
93 07 00 02 63 5C D0 10 05 05 A3 0F F5 FE E3 1D
E5 FE FD 56 63 85 0F 00 23 00 F5 01 05 05 63 08
0F 00 A1 47 63 00 F6 0E C1 47 63 03 F6 0C 19 E8
B3 07 D5 00 63 56 D0 0E 05 05 A3 0F 75 FE E3 9D
A7 FE FD 56 B3 87 08 41 AA 97 13 07 00 03 63 55
18 0D 05 05 A3 0F E5 FE E3 9D A7 FE 33 87 B2 00
3E 86 03 48 07 00 3A 85 05 06 A3 0F 06 FF 7D 17
E3 99 A2 FE 85 05 BE 95 63 5E D0 08 33 85 D5 00
93 07 00 02 85 05 A3 8F F5 FE E3 1D B5 FE 76 44
E6 44 25 61 82 80 81 4F 0D BF F9 9B A2 84 13 F8
27 00 93 03 00 02 13 FF 07 02 E3 06 08 FE 11 B7
B3 05 B0 40 FD 16 93 0F D0 02 E3 1A 0F F0 AE 87
01 48 93 02 C1 00 B3 F8 C7 02 C2 85 05 08 33 8E
02 01 3E 83 F6 98 83 C8 08 00 B3 D7 C7 02 A3 0F
1E FF E3 72 C3 FE 21 B7 FD 16 93 0F B0 02 F1 BD
93 07 00 03 23 00 F5 00 93 07 80 07 A3 00 F5 00
09 05 35 B7 93 07 00 03 23 00 F5 00 05 05 05 B7
F9 16 F1 B5 2E 85 A5 BF AA 87 89 B7 FD 16 DD BD
FD 16 0D B7
@4000451A
B7 07 00 20 C8 43 05 89 82 80
@40004524
37 07 00 20 5C 43 85 8B F5 FF 48 C7 82 80
@40004532
83 46 05 00 99 CA 37 07 00 20 05 05 5C 43 85 8B
F5 FF 54 C7 83 46 05 00 ED FA 82 80
@4000454E
37 07 00 20 5C 43 85 8B F5 FF 48 C7 82 80
@4000455C
13 01 01 B7 23 20 E1 48 23 26 11 46 23 24 81 46
23 22 91 46 23 20 21 47 23 2E 31 45 23 2C 41 45
23 2A 51 45 23 28 61 45 23 26 71 45 23 24 81 45
23 22 91 45 23 20 A1 45 23 2E B1 43 23 2A B1 46
23 2C C1 46 23 2E D1 46 23 22 F1 48 23 24 01 49
23 26 11 49 83 47 05 00 13 07 41 47 3A CA 63 8B
07 5A 93 09 01 03 2A 83 3A 8A 4E 85 13 09 50 02
C1 44 17 14 00 00 13 04 E4 50 A5 4D 93 0C E0 02
13 0D C0 04 13 0C 70 03 63 8C 27 03 23 00 F5 00
83 47 13 00 05 05 05 03 E5 FB 23 00 05 00 03 46
01 03 71 C6 CE 86 37 07 00 20 5C 43 85 8B F5 FF
50 C7 03 C6 16 00 93 87 16 00 6D C2 BE 86 F5 B7
81 47 03 46 13 00 93 05 13 00 13 07 06 FE 13 77
F7 0F 63 E7 E4 00 0A 07 22 97 18 43 22 97 02 87
13 07 06 FD 13 77 F7 0F 63 FD ED 10 13 07 A0 02
FD 56 63 0B E6 12 7D 57 63 03 96 0F 13 78 F6 0D
63 09 A8 07 13 08 F6 FB 13 78 F8 0F 63 60 0C 05
97 18 00 00 93 88 48 4B 0A 08 46 98 03 28 08 00
46 98 02 88 93 E7 17 00 2E 83 61 BF 93 E7 07 01
2E 83 41 BF 93 E7 47 00 2E 83 61 B7 93 E7 07 02
2E 83 41 B7 93 E7 87 00 2E 83 A5 BF AE 8A 93 07
50 02 63 09 F6 46 23 00 F5 00 83 C7 0A 00 05 05
63 94 07 46 23 00 05 00 03 46 01 03 05 FE 01 45
15 A8 B2 88 03 C6 15 00 93 8A 15 00 13 08 F6 FB
13 78 F8 0F E3 65 0C FD 17 13 00 00 13 03 C3 51
0A 08 1A 98 03 28 08 00 1A 98 02 88 B3 86 36 41
13 85 16 00 83 20 C1 46 03 24 81 46 83 24 41 46
03 29 01 46 83 29 C1 45 03 2A 81 45 83 2A 41 45
03 2B 01 45 83 2B C1 44 03 2C 81 44 83 2C 41 44
03 2D 01 44 83 2D C1 43 13 01 01 49 82 80 03 C6
15 00 A5 48 13 88 15 00 13 07 06 FD 13 77 F7 0F
63 F2 E8 2C 13 07 A0 02 63 03 E6 2E C2 85 01 47
F5 BD 81 46 25 48 13 97 26 00 36 97 85 05 06 07
32 97 03 C6 05 00 93 06 07 FD 13 07 06 FD 13 77
F7 0F E3 72 E8 FE C1 BD 83 26 0A 00 03 46 23 00
93 05 23 00 11 0A E3 D0 06 EC B3 06 D0 40 93 E7
07 01 55 BD 93 E7 07 04 13 07 C0 06 63 86 E8 2A
03 2E 0A 00 81 45 01 47 33 06 BE 00 03 46 06 00
3E C4 36 C6 93 0F 4A 00 93 03 30 06 97 1E 00 00
93 8E 0E 20 13 0B 40 06 A9 4B 93 02 00 03 11 43
13 0F E0 02 13 08 17 00 15 EA 93 07 07 42 18 08
3E 97 23 04 57 BE 85 05 63 83 65 08 93 07 08 42
18 08 33 86 E7 00 23 04 E6 BF 33 06 BE 00 03 46
06 00 13 07 18 00 13 08 17 00 61 DA 63 D2 C3 1C
B3 67 66 03 93 06 07 42 93 08 01 01 B6 98 C6 86
13 08 08 42 93 08 01 01 46 98 42 C2 09 07 F6 88
13 08 17 00 33 46 66 03 33 CA 77 03 76 96 03 46
06 00 23 84 C6 BE 76 9A 33 E6 77 03 03 4A 0A 00
92 47 23 84 47 BF B2 98 03 C6 08 00 93 07 07 42
18 08 3E 97 23 04 C7 BE 85 05 E3 91 65 F8 A2 47
B2 46 C1 8B 95 E3 13 86 F6 FF 63 51 D8 3A B3 87
06 41 AA 97 13 07 00 02 05 05 A3 0F E5 FE E3 9D
A7 FE B3 06 D8 40 B2 96 30 08 B3 07 05 01 2A 87
83 45 06 00 05 07 05 06 A3 0F B7 FE E3 9A E7 FE
63 57 D8 34 36 95 13 07 00 02 85 07 A3 8F E7 FE
E3 1D F5 FE 83 C7 1A 00 13 83 1A 00 7E 8A E3 95
07 D0 21 BB 93 E7 07 04 41 46 13 08 4A 00 83 25
0A 00 42 8A 9D 3C 83 C7 1A 00 13 83 1A 00 E3 95
07 CE E5 B9 AE 8A C1 8B 13 06 4A 00 13 83 1A 00
63 8F 07 22 83 27 0A 00 85 45 13 07 15 00 23 00
F5 00 93 07 00 02 36 95 63 D6 D5 30 05 07 A3 0F
F7 FE E3 1D A7 FE 83 C7 1A 00 32 8A E3 96 07 CA
6D B9 AE 8A 03 26 0A 00 11 0A 63 0D 06 1E 83 45
06 00 63 84 05 26 63 02 07 26 B2 85 29 A0 33 88
E5 40 63 07 C8 00 03 C8 15 00 85 05 E3 19 08 FE
13 F7 07 01 B3 87 C5 40 63 02 07 20 63 53 F0 2C
33 08 F6 00 2A 87 83 45 06 00 05 06 05 07 A3 0F
B7 FE E3 1A 06 FF 33 07 F5 00 33 85 F6 40 13 83
1A 00 3A 95 13 06 00 02 63 DC D7 26 05 07 A3 0F
C7 FE E3 1D A7 FE 83 C7 1A 00 E3 97 07 C2 35 B9
AE 8A 7D 56 63 8C C6 16 83 25 0A 00 41 46 11 0A
69 3A 83 C7 1A 00 13 83 1A 00 E3 97 07 C0 31 B9
A5 47 F6 88 E3 D1 C7 E8 29 4A B3 47 46 03 97 18
00 00 93 88 E8 FD 13 07 07 42 14 08 BA 96 42 87
05 08 33 66 46 03 33 8A F8 00 03 4A 0A 00 23 84
46 BF 91 BD 01 47 3A 83 13 17 23 00 1A 97 05 08
06 07 32 97 03 46 08 00 13 03 07 FD 93 05 06 FD
93 F5 F5 0F E3 F2 B8 FE 1A 87 C2 85 05 B1 03 27
0A 00 13 88 25 00 03 C6 25 00 93 45 F7 FF FD 85
6D 8F 11 0A C2 85 19 B1 13 F7 07 04 17 13 00 00
13 03 03 F7 09 C7 17 13 00 00 13 03 E3 F8 83 2E
0A 00 01 46 81 48 19 4E 13 0F A0 03 01 A8 13 87
28 42 33 08 77 00 8D 08 23 04 E8 BF 33 87 CE 00
03 47 07 00 93 03 01 01 05 06 13 58 47 00 3D 8B
1A 97 1A 98 83 4F 07 00 83 42 08 00 13 87 08 42
1E 97 23 04 57 BE A3 04 F7 BF E3 12 C6 FD C1 8B
9D E3 C5 47 13 86 F6 FF 63 D1 D7 18 93 87 F6 FE
AA 97 13 07 00 02 05 05 A3 0F E5 FE E3 1D F5 FE
15 8E 93 06 16 01 30 08 93 07 15 01 2A 87 03 48
06 00 05 07 05 06 A3 0F 07 FF E3 1A F7 FE 45 46
63 58 D6 12 36 95 13 07 00 02 85 07 A3 8F E7 FE
E3 1D F5 FE 83 C7 25 00 11 0A 13 83 25 00 E3 95
07 AC E1 BC 83 C7 0A 00 23 00 F5 00 83 C7 1A 00
05 05 13 83 1A 00 E3 99 07 AA C1 B4 93 E7 17 00
A1 46 59 B5 17 16 00 00 13 06 86 ED 29 B5 85 47
63 D4 D7 0A 93 87 F6 FF AA 97 13 07 00 02 05 05
A3 0F E5 FE E3 1D F5 FE 81 46 6D B3 93 E7 27 00
29 46 A5 BB 93 09 01 03 4E 85 41 B4 13 88 F6 FF
63 D3 D7 0C 33 87 F6 40 2A 97 93 05 00 02 05 05
A3 0F B5 FE E3 1D E5 FE B3 86 D7 40 C2 96 F9 BB
93 E7 27 00 13 08 4A 00 AE 8A 29 46 89 B3 21 46
2D BB 29 46 1D BB AE 8A E5 BE C1 8B B9 CB 2A 87
81 47 E1 BB 93 E7 07 04 AE 8A DD B6 13 08 4A 00
AE 8A 29 46 29 BB 93 E7 07 04 13 08 4A 00 AE 8A
41 46 31 B3 13 08 4A 00 AE 8A 41 46 09 B3 13 08
4A 00 AE 8A 21 46 E5 B9 83 27 0A 00 05 05 32 8A
A3 0F F5 FE 83 C7 1A 00 E3 90 07 9E FD B2 3E 85
D1 B1 13 88 F6 FF E3 47 D0 F6 13 83 1A 00 2A 87
83 C7 1A 00 3A 85 E3 91 07 9C C1 BA B2 86 AD B9
3A 85 CD B5 83 C7 1A 00 32 8A 3A 85 E3 96 07 9A
6D BA 2A 87 99 BB C2 86 15 BB B2 86 69 BD
@40004C4A
4D 71 23 24 81 14 23 20 21 15 23 2E 31 13 23 2C
41 13 23 26 11 14 23 22 91 14 23 2A 51 13 23 28
61 13 23 26 71 13 23 24 81 13 23 22 91 13 23 20
A1 13 23 2E B1 11 AA 89 2E 89 32 84 36 C6 13 0A
50 02 29 A0 31 C5 CA 85 05 04 82 99 03 45 04 00
E3 1A 45 FF 83 46 14 00 93 0A 14 00 93 07 00 02
56 87 3E C4 FD 54 7D 5B 81 45 93 87 D6 FD 93 F7
F7 0F 13 06 50 05 13 04 17 00 63 65 F6 06 17 16
00 00 13 06 86 01 8A 07 B2 97 9C 43 B2 97 82 87
83 20 C1 14 03 24 81 14 83 24 41 14 03 29 01 14
83 29 C1 13 03 2A 81 13 83 2A 41 13 03 2B 01 13
83 2B C1 12 03 2C 81 12 83 2C 41 12 03 2D 01 12
83 2D C1 11 71 61 82 80 36 C4 83 46 17 00 13 06
50 05 22 87 93 87 D6 FD 93 F7 F7 0F 13 04 17 00
E3 7F F6 F8 CA 85 13 05 50 02 82 99 56 84 B9 BF
03 46 17 00 A5 47 93 84 06 FD 13 07 06 FD B2 86
63 E8 E7 26 22 87 25 45 93 97 24 00 A6 97 05 07
86 07 B2 97 03 46 07 00 93 84 07 FD 93 07 06 FD
B2 86 E3 73 F5 FE E3 52 0B F4 26 8B FD 54 35 BF
83 46 17 00 22 87 15 BF CA 85 13 05 50 02 82 99
31 B7 B2 47 83 46 17 00 22 87 84 43 91 07 3E C6
D9 BF 13 05 00 03 CA 85 82 99 CA 85 13 05 80 07
82 99 B2 47 C1 4A 81 4D 13 87 47 00 B2 47 01 4C
84 43 3A C6 56 86 81 46 26 85 E2 85 EF D0 1F 90
2A C8 63 80 8D 1B 93 0B 41 01 85 4C 56 86 81 46
26 85 E2 85 EF D0 AF D8 56 86 81 46 AA 84 2E 8C
EF D0 DF 8D 23 A0 AB 00 66 8D 91 0B 85 0C E3 9F
8D FD E3 FD 54 FD 93 0A FB FF 93 84 FC FF 63 D8
6C 01 22 45 FD 1A CA 85 82 99 E3 9C 9A FE 93 17
2D 00 C1 07 B3 8A 27 00 A5 44 11 A0 3E 8D 03 A5
0A 00 CA 85 F1 1A B3 B7 A4 00 B3 07 F0 40 93 F7
77 02 93 87 07 03 3E 95 82 99 93 07 FD FF E3 1F
0D FC A9 B5 85 47 63 C3 B7 12 B2 47 84 43 91 07
3E C6 13 DC F4 41 63 5E 0C 00 CA 85 13 05 D0 02
82 99 33 37 90 00 B3 07 80 41 B3 04 90 40 33 8C
E7 40 A9 4A 81 4D 3D BF 83 46 17 00 85 05 22 87
2D B5 C1 4A 81 4D 85 47 63 C0 B7 0C B2 47 13 87
47 00 29 BF B2 47 83 AA 07 00 93 8B 47 00 63 8A
0A 0E 63 5D 60 07 22 47 93 07 D0 02 63 11 F7 04
03 C5 0A 00 05 C1 7D 5C 63 C5 04 00 FD 14 63 89
84 01 CA 85 85 0A 82 99 03 C5 0A 00 7D 1B 6D F5
63 59 60 01 7D 1B CA 85 13 05 00 02 82 99 E3 1B
0B FE 5E C6 65 B3 97 1A 00 00 93 8A 0A B3 D6 87
B3 86 9A 00 89 E4 29 A8 85 07 63 85 D7 00 03 C7
07 00 7D FB B3 87 57 41 33 0B FB 40 63 58 60 01
22 45 7D 1B CA 85 82 99 E3 1C 0B FE 03 C5 0A 00
69 D1 7D 5C 51 BF 93 47 FB FF FD 87 83 46 17 00
33 7B FB 00 22 87 95 BB B2 47 CA 85 88 43 93 8B
47 00 82 99 5E C6 99 B3 B2 47 93 8B 77 00 93 FB
8B FF 93 87 8B 00 83 A4 0B 00 03 AC 4B 00 3E C6
91 BD E3 F2 54 E7 01 4D 85 4C 71 B5 B2 47 93 8B
77 00 93 FB 8B FF 93 87 8B 00 83 A4 0B 00 03 AC
4B 00 3E C6 C9 BD A9 4A 81 4D F5 BD A1 4A 81 4D
DD BD 63 57 60 01 22 47 93 07 D0 02 E3 15 F7 F4
97 1A 00 00 93 8A 6A A7 13 05 80 02 7D 5C 29 B7
22 87 55 BB
@40004FBE
9C 41 23 80 A7 00 9C 41 85 07 9C C1 82 80
@40004FCC
03 28 02 04 93 07 02 00 C2 97 19 71 13 07 18 00
23 20 E2 04 23 80 A7 00 93 06 F1 03 A9 47 93 F6
06 FC 63 09 F5 00 93 07 00 04 63 05 F7 00 01 45
09 61 82 80 13 08 00 04 23 A0 06 01 81 48 23 A2
16 01 05 4E 23 A4 C6 01 81 4E 23 A6 D6 01 13 03
02 00 23 A8 66 00 81 43 23 AA 76 00 98 CE 93 58
F7 41 23 AE 16 01 0F 00 F0 0F 17 C6 FF FF 13 06
A6 FC 14 C2 81 47 5C C2 17 C6 FF FF 13 06 C6 FF
18 42 5C 42 5D 8F 6D DF 81 47 1C C2 01 48 23 22
06 01 0F 00 F0 0F 23 20 02 04 98 42 01 45 DC 42
09 61 82 80
@40005070
73 27 00 B0 97 47 00 00 93 87 87 DA 11 C5 98 C3
73 27 20 B0 D8 C3 82 80 90 43 97 46 00 00 93 86
A6 D8 11 8F 17 16 00 00 13 06 46 99 90 C2 98 C3
73 27 20 B0 D0 43 97 15 00 00 93 85 A5 98 CC C2
11 8F D8 C3 82 80
@400050B6
93 16 15 00 13 E7 16 00 97 C6 FF FF 93 86 26 F4
81 47 98 C2 DC C2 01 A0
@400050CE
05 66 97 C7 FF FF 93 87 07 F3 13 06 36 A7 81 46
90 C3 D4 C3 01 A0
@400050E4
41 11 06 C6 F9 37
@400050EA
97 C7 FF FF 93 87 67 F1 13 06 D0 10 81 46 90 C3
D4 C3 01 A0
@400050FE
83 47 05 00 19 71 13 06 F1 03 2A 88 13 76 06 FC
81 48 B5 C7 AA 87 03 C7 17 00 85 07 6D FF 33 83
A7 40 81 43 13 07 00 04 18 C2 81 47 5C C2 05 47
18 C6 81 47 5C C6 23 28 06 01 23 2A 16 01 23 2C
66 00 23 2E 76 00 0F 00 F0 0F 97 C6 FF FF 93 86
86 EB 90 C2 81 47 DC C2 97 C6 FF FF 93 86 A6 EE
98 42 DC 42 5D 8F 6D DF 81 47 9C C2 01 48 23 A2
06 01 0F 00 F0 0F 18 42 5C 42 09 61 82 80 01 43
81 43 4D B7
@40005182
01 E1 82 80
@40005186
79 71 2A 87 06 D6 68 00 93 06 B1 01 25 48 11 A0
BE 86 93 77 F7 00 B3 37 F8 00 B3 07 F0 40 93 F7
77 02 13 76 F7 00 93 87 07 03 B2 97 23 80 F6 00
13 96 C5 01 11 83 93 87 F6 FF 51 8F 91 81 E3 19
D5 FC 23 0E 01 00 0D 3F B2 50 45 61 82 80
@400051D4
39 71 13 03 41 02 2A 8E 2E D2 32 D4 36 D6 17 05
00 00 13 05 A5 DE 9A 86 72 86 81 45 06 CE 3A D8
3E DA 42 DC 46 DE 1A C6 B9 34 F2 40 01 45 21 61
82 80
@40005206
5D 71 13 03 81 03 22 D4 2A C6 32 DC 36 DE 2A 84
2E 86 17 05 00 00 13 05 65 DA 6C 00 9A 86 06 D6
BE C2 BA C0 C2 C4 C6 C6 1A CE 29 3C B2 47 23 80
07 00 32 45 B2 50 01 8D 22 54 61 61 82 80
@40005244
B3 67 B5 00 D1 8F 8D 8B B3 06 C5 00 91 CF 2E 96
AA 87 63 76 D5 02 03 C7 05 00 85 05 85 07 A3 8F
E7 FE E3 1A B6 FE 82 80 E3 7F D5 FE AA 87 98 41
91 07 91 05 23 AE E7 FE E3 EB D7 FE 82 80 82 80
@40005284
B3 67 C5 00 8D 8B 2A 96 81 CF 93 F5 F5 0F AA 87
63 79 C5 02 85 07 A3 8F B7 FE E3 9D C7 FE 82 80
93 F5 F5 0F 13 97 85 00 2E 97 93 17 07 01 3E 97
E3 77 C5 FE AA 87 91 07 23 AE E7 FE E3 ED C7 FE
82 80 82 80
@400052C8
35 71 97 47 00 00 93 87 A7 B5 52 C5 17 4A 00 00
13 0A 0A B5 4E C7 B3 09 FA 40 26 CB 4A C9 AA 84
2E 89 12 85 BE 85 4E 86 06 CF 22 CD 56 C3 92 8A
B1 37 13 86 C1 89 33 06 46 41 81 45 33 85 3A 01
B5 3F CA 85 26 85 95 3D 81 45 01 45 EF D0 9F D2
17 49 00 00 13 09 49 B0 83 26 09 00 13 04 F1 03
13 74 04 FC AA 84 8D EA 83 26 49 00 99 E2 26 85
BD 3B 22 89 97 49 00 00 93 89 89 AD 03 A6 49 00
4A 85 97 05 00 00 93 85 A5 70 55 3D 2A 99 E3 00
24 FF 22 85 4D 33 E1 BF 97 49 00 00 93 89 49 AB
03 A6 09 00 97 05 00 00 93 85 85 6E 22 85 41 3D
83 26 49 00 33 09 A4 00 F9 DA C9 B7
@40005384
83 47 05 00 89 CB AA 87 03 C7 17 00 85 07 6D FF
33 85 A7 40 82 80 01 45 82 80
@4000539E
B3 06 B5 00 AA 87 89 E5 29 A8 85 07 63 88 F6 00
03 C7 07 00 7D FB 33 85 A7 40 82 80 33 85 A6 40
82 80 01 45 82 80
@400053C4
83 47 05 00 85 05 05 05 03 C7 F5 FF 91 C7 E3 89
E7 FE 33 85 E7 40 82 80 81 47 E5 BF
@400053E0
AA 87 03 C7 05 00 85 07 85 05 A3 8F E7 FE 75 FB
82 80
@400053F2
03 47 05 00 93 06 00 02 AA 87 63 17 D7 00 03 C7
17 00 85 07 E3 0D D7 FE 93 06 D0 02 63 02 D7 04
93 06 B0 02 63 07 D7 02 83 C6 07 00 81 45 9D C6
01 45 85 07 13 17 25 00 13 86 06 FD 83 C6 07 00
2A 97 06 07 33 05 E6 00 ED F6 91 C9 33 05 A0 40
82 80 83 C6 17 00 81 45 85 07 F9 FA 01 45 82 80
83 C6 17 00 85 45 85 07 E1 F6 01 45 CD BF
@40005460
70 69 6B 61 63 68 75 0A 00 00 00 00 36 6B 20 70
65 72 66 6F 72 6D 61 6E 63 65 20 72 75 6E 20 70
61 72 61 6D 65 74 65 72 73 20 66 6F 72 20 63 6F
72 65 6D 61 72 6B 2E 0A 00 00 00 00 36 6B 20 76
61 6C 69 64 61 74 69 6F 6E 20 72 75 6E 20 70 61
72 61 6D 65 74 65 72 73 20 66 6F 72 20 63 6F 72
65 6D 61 72 6B 2E 0A 00 50 72 6F 66 69 6C 65 20
67 65 6E 65 72 61 74 69 6F 6E 20 72 75 6E 20 70
61 72 61 6D 65 74 65 72 73 20 66 6F 72 20 63 6F
72 65 6D 61 72 6B 2E 0A 00 00 00 00 32 4B 20 70
65 72 66 6F 72 6D 61 6E 63 65 20 72 75 6E 20 70
61 72 61 6D 65 74 65 72 73 20 66 6F 72 20 63 6F
72 65 6D 61 72 6B 2E 0A 00 00 00 00 32 4B 20 76
61 6C 69 64 61 74 69 6F 6E 20 72 75 6E 20 70 61
72 61 6D 65 74 65 72 73 20 66 6F 72 20 63 6F 72
65 6D 61 72 6B 2E 0A 00 5B 25 75 5D 45 52 52 4F
52 21 20 6C 69 73 74 20 63 72 63 20 30 78 25 30
34 78 20 2D 20 73 68 6F 75 6C 64 20 62 65 20 30
78 25 30 34 78 0A 00 00 5B 25 75 5D 45 52 52 4F
52 21 20 6D 61 74 72 69 78 20 63 72 63 20 30 78
25 30 34 78 20 2D 20 73 68 6F 75 6C 64 20 62 65
20 30 78 25 30 34 78 0A 00 00 00 00 5B 25 75 5D
45 52 52 4F 52 21 20 73 74 61 74 65 20 63 72 63
20 30 78 25 30 34 78 20 2D 20 73 68 6F 75 6C 64
20 62 65 20 30 78 25 30 34 78 0A 00 43 6F 72 65
4D 61 72 6B 20 53 69 7A 65 20 20 20 20 3A 20 25
6C 75 0A 00 54 6F 74 61 6C 20 74 69 63 6B 73 20
20 20 20 20 20 3A 20 25 4C 75 0A 00 54 6F 74 61
6C 20 74 69 6D 65 20 28 73 65 63 73 29 3A 20 25
64 0A 00 00 49 74 65 72 61 74 69 6F 6E 73 2F 53
65 63 20 20 20 3A 20 25 64 0A 00 00 45 52 52 4F
52 21 20 4D 75 73 74 20 65 78 65 63 75 74 65 20
66 6F 72 20 61 74 20 6C 65 61 73 74 20 31 30 20
73 65 63 73 20 66 6F 72 20 61 20 76 61 6C 69 64
20 72 65 73 75 6C 74 21 0A 00 00 00 49 74 65 72
61 74 69 6F 6E 73 20 20 20 20 20 20 20 3A 20 25
6C 75 0A 00 47 43 43 31 32 2E 32 2E 30 00 00 00
43 6F 6D 70 69 6C 65 72 20 76 65 72 73 69 6F 6E
20 3A 20 25 73 0A 00 00 2D 4F 32 20 2D 6D 63 6D
6F 64 65 6C 3D 6D 65 64 61 6E 79 20 2D 73 74 61
74 69 63 20 2D 73 74 64 3D 67 6E 75 39 39 20 2D
66 6E 6F 2D 63 6F 6D 6D 6F 6E 20 2D 6E 6F 73 74
64 6C 69 62 20 2D 6E 6F 73 74 61 72 74 66 69 6C
65 73 20 2D 66 6E 6F 2D 62 75 69 6C 74 69 6E 20
2D 66 66 75 6E 63 74 69 6F 6E 2D 73 65 63 74 69
6F 6E 73 20 2D 6C 6D 20 2D 6C 67 63 63 20 2D 54
20 72 69 73 63 76 33 32 2D 62 61 72 65 6D 65 74
61 6C 2F 6C 69 6E 6B 64 65 6E 65 2E 6C 64 20 2D
44 50 45 52 46 4F 52 4D 41 4E 43 45 5F 52 55 4E
3D 31 20 20 00 00 00 00 43 6F 6D 70 69 6C 65 72
20 66 6C 61 67 73 20 20 20 3A 20 25 73 0A 00 00
53 54 41 43 4B 00 00 00 4D 65 6D 6F 72 79 20 6C
6F 63 61 74 69 6F 6E 20 20 3A 20 25 73 0A 00 00
73 65 65 64 63 72 63 20 20 20 20 20 20 20 20 20
20 3A 20 30 78 25 30 34 78 0A 00 00 5B 25 64 5D
63 72 63 6C 69 73 74 20 20 20 20 20 20 20 3A 20
30 78 25 30 34 78 0A 00 5B 25 64 5D 63 72 63 6D
61 74 72 69 78 20 20 20 20 20 3A 20 30 78 25 30
34 78 0A 00 5B 25 64 5D 63 72 63 73 74 61 74 65
20 20 20 20 20 20 3A 20 30 78 25 30 34 78 0A 00
5B 25 64 5D 63 72 63 66 69 6E 61 6C 20 20 20 20
20 20 3A 20 30 78 25 30 34 78 0A 00 43 6F 72 72
65 63 74 20 6F 70 65 72 61 74 69 6F 6E 20 76 61
6C 69 64 61 74 65 64 2E 20 53 65 65 20 52 45 41
44 4D 45 2E 6D 64 20 66 6F 72 20 72 75 6E 20 61
6E 64 20 72 65 70 6F 72 74 69 6E 67 20 72 75 6C
65 73 2E 0A 00 00 00 00 43 61 6E 6E 6F 74 20 76
61 6C 69 64 61 74 65 20 6F 70 65 72 61 74 69 6F
6E 20 66 6F 72 20 74 68 65 73 65 20 73 65 65 64
20 76 61 6C 75 65 73 2C 20 70 6C 65 61 73 65 20
63 6F 6D 70 61 72 65 20 77 69 74 68 20 72 65 73
75 6C 74 73 20 6F 6E 20 61 20 6B 6E 6F 77 6E 20
70 6C 61 74 66 6F 72 6D 2E 0A 00 00 45 72 72 6F
72 73 20 64 65 74 65 63 74 65 64 0A 00 00 00 00
53 74 61 74 69 63 00 00 48 65 61 70 00 00 00 00
53 74 61 63 6B 00 00 00 54 30 2E 33 65 2D 31 46
00 00 00 00 2D 54 2E 54 2B 2B 54 71 00 00 00 00
31 54 33 2E 34 65 34 7A 00 00 00 00 33 34 2E 30
65 2D 54 5E 00 00 00 00 35 2E 35 30 30 65 2B 33
00 00 00 00 2D 2E 31 32 33 65 2D 32 00 00 00 00
2D 38 37 65 2B 38 33 32 00 00 00 00 2B 30 2E 36
65 2D 31 32 00 00 00 00 33 35 2E 35 34 34 30 30
00 00 00 00 2E 31 32 33 34 35 30 30 00 00 00 00
2D 31 31 30 2E 37 30 30 00 00 00 00 2B 30 2E 36
34 34 30 30 00 00 00 00 35 30 31 32 00 00 00 00
31 32 33 34 00 00 00 00 2D 38 37 34 00 00 00 00
2B 31 32 32 00 00 00 00 30 31 32 33 34 35 36 37
38 39 61 62 63 64 65 66 67 68 69 6A 6B 6C 6D 6E
6F 70 71 72 73 74 75 76 77 78 79 7A 00 00 00 00
30 31 32 33 34 35 36 37 38 39 41 42 43 44 45 46
47 48 49 4A 4B 4C 4D 4E 4F 50 51 52 53 54 55 56
57 58 59 5A 00 00 00 00 3C 4E 55 4C 4C 3E 00 00
28 6E 75 6C 6C 29 00 00 6D 63 79 63 6C 65 00 00
6D 69 6E 73 74 72 65 74 00 00 00 00 49 6D 70 6C
65 6D 65 6E 74 20 6D 61 69 6E 28 29 2C 20 66 6F
6F 21 0A 00 25 73 20 3D 20 25 64 0A 00
@40005A60
B0 D4 40 33 79 6A 14 E7 C1 E3 00 00 52 BE 99 11
08 56 D7 1F 47 07 00 00 47 5E BF 39 A4 E5 3A 8E
84 8D 00 00 A8 59 00 40 B0 59 00 40 B8 59 00 40
C0 59 00 40 78 59 00 40 84 59 00 40 90 59 00 40
9C 59 00 40 48 59 00 40 54 59 00 40 60 59 00 40
6C 59 00 40 18 59 00 40 24 59 00 40 30 59 00 40
3C 59 00 40 66 E6 FF FF 42 E6 FF FF 4C E6 FF FF
56 E6 FF FF 5C E6 FF FF 38 E6 FF FF C4 EB FF FF
60 EB FF FF 60 EB FF FF BC EB FF FF 60 EB FF FF
60 EB FF FF 60 EB FF FF 60 EB FF FF 60 EB FF FF
60 EB FF FF 60 EB FF FF B4 EB FF FF 60 EB FF FF
AC EB FF FF 60 EB FF FF 60 EB FF FF A4 EB FF FF
A0 F0 FF FF 88 EB FF FF 88 EB FF FF 88 EB FF FF
88 EB FF FF 88 EB FF FF 88 EB FF FF 88 EB FF FF
88 EB FF FF 88 EB FF FF 88 EB FF FF 88 EB FF FF
88 EB FF FF 88 EB FF FF 88 EB FF FF 88 EB FF FF
88 EB FF FF 88 EB FF FF 88 EB FF FF 88 EB FF FF
88 EB FF FF 88 EB FF FF 88 EB FF FF B2 F0 FF FF
88 EB FF FF 88 EB FF FF 88 EB FF FF 88 EB FF FF
88 EB FF FF 88 EB FF FF 88 EB FF FF 88 EB FF FF
92 F0 FF FF 88 EB FF FF E0 ED FF FF 7C F0 FF FF
88 EB FF FF 88 EB FF FF 88 EB FF FF 88 EB FF FF
7C F0 FF FF 88 EB FF FF 88 EB FF FF 88 EB FF FF
88 EB FF FF 88 EB FF FF CA F0 FF FF 9C EE FF FF
88 EB FF FF 88 EB FF FF 1E EE FF FF 88 EB FF FF
A8 F0 FF FF 88 EB FF FF 88 EB FF FF C0 F0 FF FF
A0 EB FF FF AA EA FF FF AA EA FF FF AA EA FF FF
AA EA FF FF AA EA FF FF AA EA FF FF AA EA FF FF
AA EA FF FF AA EA FF FF AA EA FF FF AA EA FF FF
AA EA FF FF AA EA FF FF AA EA FF FF AA EA FF FF
AA EA FF FF AA EA FF FF AA EA FF FF AA EA FF FF
AA EA FF FF AA EA FF FF AA EA FF FF E0 EC FF FF
AA EA FF FF AA EA FF FF AA EA FF FF AA EA FF FF
AA EA FF FF AA EA FF FF AA EA FF FF AA EA FF FF
A4 EB FF FF AA EA FF FF 02 ED FF FF 68 EF FF FF
AA EA FF FF AA EA FF FF AA EA FF FF AA EA FF FF
68 EF FF FF AA EA FF FF AA EA FF FF AA EA FF FF
AA EA FF FF AA EA FF FF AA EF FF FF BE ED FF FF
AA EA FF FF AA EA FF FF 40 ED FF FF AA EA FF FF
AE EF FF FF AA EA FF FF AA EA FF FF E4 EC FF FF
9A F0 FF FF 4E F0 FF FF A2 F0 FF FF 4E F0 FF FF
4E F0 FF FF 4E F0 FF FF 4E F0 FF FF AC F0 FF FF
4E F0 FF FF 4E F0 FF FF 32 F0 FF FF 50 F2 FF FF
4E F0 FF FF 32 F0 FF FF 5A F0 FF FF 5A F0 FF FF
5A F0 FF FF 5A F0 FF FF 5A F0 FF FF 5A F0 FF FF
5A F0 FF FF 5A F0 FF FF 5A F0 FF FF 4E F0 FF FF
4E F0 FF FF 4E F0 FF FF 4E F0 FF FF 4E F0 FF FF
4E F0 FF FF 4E F0 FF FF 4E F0 FF FF 4E F0 FF FF
4E F0 FF FF 4E F0 FF FF 4E F0 FF FF 4E F0 FF FF
4E F0 FF FF 4E F0 FF FF 4E F0 FF FF 4E F0 FF FF
4E F0 FF FF 4E F0 FF FF 4E F0 FF FF 4E F0 FF FF
4E F0 FF FF 4E F0 FF FF 4E F0 FF FF 4E F0 FF FF
4E F0 FF FF 4E F0 FF FF 4E F0 FF FF 4E F0 FF FF
4E F0 FF FF 4E F0 FF FF 4E F0 FF FF 4E F0 FF FF
4E F0 FF FF 4E F0 FF FF 4E F0 FF FF 4E F0 FF FF
4E F0 FF FF 4E F0 FF FF 4E F0 FF FF 4E F0 FF FF
62 F2 FF FF 6E F1 FF FF 4E F0 FF FF 4E F0 FF FF
4E F0 FF FF 4E F0 FF FF 4E F0 FF FF 4E F0 FF FF
4E F0 FF FF A2 F1 FF FF 4E F0 FF FF 4E F0 FF FF
B6 F2 FF FF BC F0 FF FF 4E F0 FF FF 4E F0 FF FF
BE F1 FF FF 4E F0 FF FF B0 F2 FF FF 4E F0 FF FF
4E F0 FF FF AC F1 FF FF 00 01 02 02 03 03 03 03
04 04 04 04 04 04 04 04 05 05 05 05 05 05 05 05
05 05 05 05 05 05 05 05 06 06 06 06 06 06 06 06
06 06 06 06 06 06 06 06 06 06 06 06 06 06 06 06
06 06 06 06 06 06 06 06 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07
07 07 07 07 07 07 07 07 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08 08 08 08 08 08 08 08 08
08 08 08 08 08 08 08 08
@40005F38
10 00 00 00 00 00 00 00 03 7A 52 00 01 7C 01 01
1B 0D 02 00 10 00 00 00 18 00 00 00 AC C0 FF FF
68 03 00 00 00 00 00 00 10 00 00 00 2C 00 00 00
00 C4 FF FF 5E 03 00 00 00 00 00 00 10 00 00 00
40 00 00 00 4A C7 FF FF 28 03 00 00 00 00 00 00
@40005F88
00 59 00 40 08 59 00 40 10 59 00 40 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 0A 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 0A 20 20
20 20 20 20 20 20 20 20 20 20 20 20 4F 4F 4F 4F
4F 4F 4F 4F 4F 20 20 20 20 20 20 20 20 20 20 20
20 20 47 47 47 47 47 47 47 47 47 47 47 47 47 55
55 55 55 55 55 55 55 20 20 20 20 20 55 55 55 55
55 55 55 55 5A 5A 5A 5A 5A 5A 5A 5A 5A 5A 5A 5A
5A 5A 5A 5A 5A 5A 5A 20 20 20 20 20 45 45 45 45
45 45 45 45 45 45 45 45 45 45 45 45 45 45 45 45
45 45 52 52 52 52 52 52 52 52 52 52 52 52 52 52
52 52 52 20 20 20 20 20 20 20 20 20 20 20 47 47
47 47 47 47 47 47 47 47 47 47 47 49 49 49 49 49
49 49 49 49 49 4E 4E 4E 4E 4E 4E 4E 4E 20 20 20
20 20 20 20 20 4E 4E 4E 4E 4E 4E 4E 4E 20 20 20
20 20 20 20 20 20 0A 20 20 20 20 20 20 20 20 20
20 20 20 4F 4F 3A 3A 3A 3A 3A 3A 3A 3A 3A 4F 4F
20 20 20 20 20 20 20 20 47 47 47 3A 3A 3A 3A 3A
3A 3A 3A 3A 3A 3A 3A 47 55 3A 3A 3A 3A 3A 3A 55
20 20 20 20 20 55 3A 3A 3A 3A 3A 3A 55 5A 3A 3A
3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 5A
20 20 20 20 20 45 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A
3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 45 52 3A 3A 3A 3A
3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 52 20 20 20
20 20 20 20 47 47 47 3A 3A 3A 3A 3A 3A 3A 3A 3A
3A 3A 3A 47 49 3A 3A 3A 3A 3A 3A 3A 3A 49 4E 3A
3A 3A 3A 3A 3A 3A 4E 20 20 20 20 20 20 20 4E 3A
3A 3A 3A 3A 3A 4E 20 20 20 20 20 20 20 20 20 0A
20 20 20 20 20 20 20 20 20 20 4F 4F 3A 3A 3A 3A
3A 3A 3A 3A 3A 3A 3A 3A 3A 4F 4F 20 20 20 20 47
47 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A
47 55 3A 3A 3A 3A 3A 3A 55 20 20 20 20 20 55 3A
3A 3A 3A 3A 3A 55 5A 3A 3A 3A 3A 3A 3A 3A 3A 3A
3A 3A 3A 3A 3A 3A 3A 3A 5A 20 20 20 20 20 45 3A
3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A
3A 3A 3A 45 52 3A 3A 3A 3A 3A 3A 52 52 52 52 52
52 3A 3A 3A 3A 3A 52 20 20 20 20 47 47 3A 3A 3A
3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 47 49 3A 3A
3A 3A 3A 3A 3A 3A 49 4E 3A 3A 3A 3A 3A 3A 3A 3A
4E 20 20 20 20 20 20 4E 3A 3A 3A 3A 3A 3A 4E 20
20 20 20 20 20 20 20 20 0A 20 20 20 20 20 20 20
20 20 4F 3A 3A 3A 3A 3A 3A 3A 4F 4F 4F 3A 3A 3A
3A 3A 3A 3A 4F 20 20 47 3A 3A 3A 3A 3A 47 47 47
47 47 47 47 47 3A 3A 3A 3A 47 55 55 3A 3A 3A 3A
3A 55 20 20 20 20 20 55 3A 3A 3A 3A 3A 55 55 5A
3A 3A 3A 5A 5A 5A 5A 5A 5A 5A 5A 3A 3A 3A 3A 3A
5A 20 20 20 20 20 20 45 45 3A 3A 3A 3A 3A 3A 45
45 45 45 45 45 45 45 45 3A 3A 3A 3A 45 52 52 3A
3A 3A 3A 3A 52 20 20 20 20 20 52 3A 3A 3A 3A 3A
52 20 20 47 3A 3A 3A 3A 3A 47 47 47 47 47 47 47
47 3A 3A 3A 3A 47 49 49 3A 3A 3A 3A 3A 3A 49 49
4E 3A 3A 3A 3A 3A 3A 3A 3A 3A 4E 20 20 20 20 20
4E 3A 3A 3A 3A 3A 3A 4E 20 20 20 20 20 20 20 20
20 0A 20 20 20 20 20 20 20 20 20 4F 3A 3A 3A 3A
3A 3A 4F 20 20 20 4F 3A 3A 3A 3A 3A 3A 4F 20 47
3A 3A 3A 3A 3A 47 20 20 20 20 20 20 20 47 47 47
47 47 47 20 55 3A 3A 3A 3A 3A 55 20 20 20 20 20
55 3A 3A 3A 3A 3A 55 20 5A 5A 5A 5A 5A 20 20 20
20 20 5A 3A 3A 3A 3A 3A 5A 20 20 20 20 20 20 20
20 20 45 3A 3A 3A 3A 3A 45 20 20 20 20 20 20 20
45 45 45 45 45 45 20 20 52 3A 3A 3A 3A 52 20 20
20 20 20 52 3A 3A 3A 3A 3A 52 20 47 3A 3A 3A 3A
3A 47 20 20 20 20 20 20 20 47 47 47 47 47 47 20
20 49 3A 3A 3A 3A 49 20 20 4E 3A 3A 3A 3A 3A 3A
3A 3A 3A 3A 4E 20 20 20 20 4E 3A 3A 3A 3A 3A 3A
4E 20 20 20 20 20 20 20 20 20 0A 20 20 20 20 20
20 20 20 20 4F 3A 3A 3A 3A 3A 4F 20 20 20 20 20
4F 3A 3A 3A 3A 3A 4F 47 3A 3A 3A 3A 3A 47 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 55 3A 3A
3A 3A 3A 44 20 20 20 20 20 44 3A 3A 3A 3A 3A 55
20 20 20 20 20 20 20 20 20 5A 3A 3A 3A 3A 3A 5A
20 20 20 20 20 20 20 20 20 20 20 45 3A 3A 3A 3A
3A 45 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 52 3A 3A 3A 3A 52 20 20 20 20 20 52 3A 3A 3A
3A 3A 52 47 3A 3A 3A 3A 3A 47 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 49 3A 3A 3A 3A 49
20 20 4E 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 4E 20
20 20 4E 3A 3A 3A 3A 3A 3A 4E 20 20 20 20 20 20
20 20 20 0A 20 20 20 20 20 20 20 20 20 4F 3A 3A
3A 3A 3A 4F 20 20 20 20 20 4F 3A 3A 3A 3A 3A 4F
47 3A 3A 3A 3A 3A 47 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 55 3A 3A 3A 3A 3A 44 20 20 20
20 20 44 3A 3A 3A 3A 3A 55 20 20 20 20 20 20 20
20 5A 3A 3A 3A 3A 3A 5A 20 20 20 20 20 20 20 20
20 20 20 20 45 3A 3A 3A 3A 3A 3A 45 45 45 45 45
45 45 45 45 45 20 20 20 20 20 52 3A 3A 3A 3A 52
52 52 52 52 52 3A 3A 3A 3A 3A 52 20 47 3A 3A 3A
3A 3A 47 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 49 3A 3A 3A 3A 49 20 20 4E 3A 3A 3A 3A
3A 3A 3A 4E 3A 3A 3A 3A 4E 20 20 4E 3A 3A 3A 3A
3A 3A 4E 20 20 20 20 20 20 20 20 20 0A 20 20 20
20 20 20 20 20 20 4F 3A 3A 3A 3A 3A 4F 20 20 20
20 20 4F 3A 3A 3A 3A 3A 4F 47 3A 3A 3A 3A 3A 47
20 20 20 20 47 47 47 47 47 47 47 47 47 47 20 55
3A 3A 3A 3A 3A 44 20 20 20 20 20 44 3A 3A 3A 3A
3A 55 20 20 20 20 20 20 20 5A 3A 3A 3A 3A 3A 5A
20 20 20 20 20 20 20 20 20 20 20 20 20 45 3A 3A
3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 45 20 20
20 20 20 52 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A
3A 52 52 20 20 47 3A 3A 3A 3A 3A 47 20 20 20 20
47 47 47 47 47 47 47 47 47 47 20 20 49 3A 3A 3A
3A 49 20 20 4E 3A 3A 3A 3A 3A 3A 4E 20 4E 3A 3A
3A 3A 4E 20 4E 3A 3A 3A 3A 3A 3A 4E 20 20 20 20
20 20 20 20 20 0A 20 20 20 20 20 20 20 20 20 4F
3A 3A 3A 3A 3A 4F 20 20 20 20 20 4F 3A 3A 3A 3A
3A 4F 47 3A 3A 3A 3A 3A 47 20 20 20 20 47 3A 3A
3A 3A 3A 3A 3A 3A 47 20 55 3A 3A 3A 3A 3A 44 20
20 20 20 20 44 3A 3A 3A 3A 3A 55 20 20 20 20 20
20 5A 3A 3A 3A 3A 3A 5A 20 20 20 20 20 20 20 20
20 20 20 20 20 20 45 3A 3A 3A 3A 3A 3A 3A 3A 3A
3A 3A 3A 3A 3A 3A 45 20 20 20 20 20 52 3A 3A 3A
3A 52 52 52 52 52 52 3A 3A 3A 3A 3A 52 20 47 3A
3A 3A 3A 3A 47 20 20 20 20 47 3A 3A 3A 3A 3A 3A
3A 3A 47 20 20 49 3A 3A 3A 3A 49 20 20 4E 3A 3A
3A 3A 3A 3A 4E 20 20 4E 3A 3A 3A 3A 4E 3A 3A 3A
3A 3A 3A 3A 4E 20 20 20 20 20 20 20 20 20 0A 20
20 20 20 20 20 20 20 20 4F 3A 3A 3A 3A 3A 4F 20
20 20 20 20 4F 3A 3A 3A 3A 3A 4F 47 3A 3A 3A 3A
3A 47 20 20 20 20 47 47 47 47 47 3A 3A 3A 3A 47
20 55 3A 3A 3A 3A 3A 44 20 20 20 20 20 44 3A 3A
3A 3A 3A 55 20 20 20 20 20 5A 3A 3A 3A 3A 3A 5A
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 45
3A 3A 3A 3A 3A 3A 45 45 45 45 45 45 45 45 45 45
20 20 20 20 20 52 3A 3A 3A 3A 52 20 20 20 20 20
52 3A 3A 3A 3A 3A 52 47 3A 3A 3A 3A 3A 47 20 20
20 20 47 47 47 47 47 3A 3A 3A 3A 47 20 20 49 3A
3A 3A 3A 49 20 20 4E 3A 3A 3A 3A 3A 3A 4E 20 20
20 4E 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 4E 20 20
20 20 20 20 20 20 20 0A 20 20 20 20 20 20 20 20
20 4F 3A 3A 3A 3A 3A 4F 20 20 20 20 20 4F 3A 3A
3A 3A 3A 4F 47 3A 3A 3A 3A 3A 47 20 20 20 20 20
20 20 20 47 3A 3A 3A 3A 47 20 55 3A 3A 3A 3A 3A
44 20 20 20 20 20 44 3A 3A 3A 3A 3A 55 20 20 20
20 5A 3A 3A 3A 3A 3A 5A 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 45 3A 3A 3A 3A 3A 45 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 52 3A
3A 3A 3A 52 20 20 20 20 20 52 3A 3A 3A 3A 3A 52
47 3A 3A 3A 3A 3A 47 20 20 20 20 20 20 20 20 47
3A 3A 3A 3A 47 20 20 49 3A 3A 3A 3A 49 20 20 4E
3A 3A 3A 3A 3A 3A 4E 20 20 20 20 4E 3A 3A 3A 3A
3A 3A 3A 3A 3A 3A 4E 20 20 20 20 20 20 20 20 20
0A 20 20 20 20 20 20 20 20 20 4F 3A 3A 3A 3A 3A
3A 4F 20 20 20 4F 3A 3A 3A 3A 3A 3A 4F 20 47 3A
3A 3A 3A 3A 47 20 20 20 20 20 20 20 47 3A 3A 3A
3A 47 20 55 3A 3A 3A 3A 3A 3A 55 20 20 20 55 3A
3A 3A 3A 3A 3A 55 20 5A 5A 5A 3A 3A 3A 3A 3A 5A
20 20 20 20 20 5A 5A 5A 5A 5A 20 20 20 20 20 20
20 45 3A 3A 3A 3A 3A 45 20 20 20 20 20 20 20 45
45 45 45 45 45 20 20 52 3A 3A 3A 3A 52 20 20 20
20 20 52 3A 3A 3A 3A 3A 52 20 47 3A 3A 3A 3A 3A
47 20 20 20 20 20 20 20 47 3A 3A 3A 3A 47 20 20
49 3A 3A 3A 3A 49 20 20 4E 3A 3A 3A 3A 3A 3A 4E
20 20 20 20 20 4E 3A 3A 3A 3A 3A 3A 3A 3A 3A 4E
20 20 20 20 20 20 20 20 20 0A 20 20 20 20 20 20
20 20 20 4F 3A 3A 3A 3A 3A 3A 3A 4F 4F 4F 3A 3A
3A 3A 3A 3A 3A 4F 20 20 47 3A 3A 3A 3A 3A 47 47
47 47 47 47 47 47 3A 3A 3A 3A 47 20 55 3A 3A 3A
3A 3A 3A 3A 55 55 55 3A 3A 3A 3A 3A 3A 3A 55 20
5A 3A 3A 3A 3A 3A 3A 5A 5A 5A 5A 5A 5A 5A 5A 3A
3A 3A 5A 20 20 20 20 20 45 45 3A 3A 3A 3A 3A 3A
45 45 45 45 45 45 45 45 3A 3A 3A 3A 3A 45 52 52
3A 3A 3A 3A 3A 52 20 20 20 20 20 52 3A 3A 3A 3A
3A 52 20 20 47 3A 3A 3A 3A 3A 47 47 47 47 47 47
47 47 3A 3A 3A 3A 47 49 49 3A 3A 3A 3A 3A 3A 49
49 4E 3A 3A 3A 3A 3A 3A 4E 20 20 20 20 20 20 4E
3A 3A 3A 3A 3A 3A 3A 3A 4E 20 20 20 20 20 20 20
20 20 0A 20 20 20 20 20 20 20 20 20 20 4F 4F 3A
3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 4F 4F 20 20
20 20 47 47 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A
3A 3A 3A 47 20 20 55 55 3A 3A 3A 3A 3A 3A 3A 3A
3A 3A 3A 3A 3A 55 55 20 20 5A 3A 3A 3A 3A 3A 3A
3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 5A 20 20 20 20
20 45 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A
3A 3A 3A 3A 3A 3A 45 52 3A 3A 3A 3A 3A 3A 52 20
20 20 20 20 52 3A 3A 3A 3A 3A 52 20 20 20 47 47
3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 47
49 3A 3A 3A 3A 3A 3A 3A 3A 49 4E 3A 3A 3A 3A 3A
3A 4E 20 20 20 20 20 20 20 4E 3A 3A 3A 3A 3A 3A
3A 4E 20 20 20 20 20 20 20 20 20 0A 20 20 20 20
20 20 20 20 20 20 20 20 4F 4F 3A 3A 3A 3A 3A 3A
3A 3A 3A 4F 4F 20 20 20 20 20 20 20 20 47 47 47
3A 3A 3A 3A 3A 3A 47 47 47 3A 3A 3A 47 20 20 20
20 55 55 3A 3A 3A 3A 3A 3A 3A 3A 3A 55 55 20 20
20 20 5A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A
3A 3A 3A 3A 5A 20 20 20 20 20 45 3A 3A 3A 3A 3A
3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 3A 45
52 3A 3A 3A 3A 3A 3A 52 20 20 20 20 20 52 3A 3A
3A 3A 3A 52 20 20 20 20 20 47 47 47 3A 3A 3A 3A
3A 3A 47 47 47 3A 3A 3A 47 49 3A 3A 3A 3A 3A 3A
3A 3A 49 4E 3A 3A 3A 3A 3A 3A 4E 20 20 20 20 20
20 20 20 4E 3A 3A 3A 3A 3A 3A 4E 20 20 20 20 20
20 20 20 20 0A 20 20 20 20 20 20 20 20 20 20 20
20 20 20 4F 4F 4F 4F 4F 4F 4F 4F 4F 20 20 20 20
20 20 20 20 20 20 20 20 20 47 47 47 47 47 47 20
20 20 47 47 47 47 20 20 20 20 20 20 55 55 55 55
55 55 55 55 55 20 20 20 20 20 20 5A 5A 5A 5A 5A
5A 5A 5A 5A 5A 5A 5A 5A 5A 5A 5A 5A 5A 5A 20 20
20 20 20 45 45 45 45 45 45 45 45 45 45 45 45 45
45 45 45 45 45 45 45 45 45 52 52 52 52 52 52 52
52 20 20 20 20 20 52 52 52 52 52 52 52 20 20 20
20 20 20 20 20 47 47 47 47 47 47 20 20 20 47 47
47 47 49 49 49 49 49 49 49 49 49 49 4E 4E 4E 4E
4E 4E 4E 4E 20 20 20 20 20 20 20 20 20 4E 4E 4E
4E 4E 4E 4E 20 20 20 20 20 20 20 20 20 0A 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 0A 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 2E 2A 2E 2C 2E 2F 2C 2C 2E 2F 2A
2C 2A 2A 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 0A
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 2C 2A 28 2F 2A
2C 23 23 23 23 23 25 25 25 25 25 26 26 26 26 25
23 23 2A 2E 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 0A 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 28 25 25 25 26 26 25 28 2A 2A 2A 2A 2A 2A 2A
2A 2A 2A 2A 2A 2A 2F 2F 23 25 25 25 25 25 28 23
2C 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 0A 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 2F 26 26 26 28 2A 2A 2A 2C
2C 2C 2C 2C 2A 2C 2A 2C 2C 2C 2C 2C 2C 2C 2C 2C
2C 2C 2C 2C 2C 2A 2F 25 25 25 25 2C 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 0A 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 2A 26 25
2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C
2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C
2C 2C 2A 28 25 23 23 25 2C 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 0A 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 2E 2C 2A 2F 2F 2F 2F 2F 2F 2A 2C
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 2C 25 25 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C
2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2E 2E 2E 2E 2E 2E
2C 2E 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 28 25
26 23 23 25 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 0A 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 2E 28 23 25 25 25 25 25 25 23 23 23 23
28 28 28 28 23 23 23 23 25 25 25 25 25 25 25 23
2A 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 23 28 2C 2C 2C
2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C
2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2C 2E 2E 2C
2C 2C 2C 2C 2E 2C 2C 2C 2A 28 26 26 25 26 28 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 0A 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 2C 23 25 25 25 23 2A 2E 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 2C 23 25 25 25 25 2C 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 2F 28 2A 2A 2A 2C 2C 2C 2C 2C 2C 2C 2C 2C
2C 2C 2C 2C 2C 2E 2C 2C 2C 2E 2E 2E 2E 2E 2E 2E
2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2C 2E 2E 2C 2C
2C 2C 2C 2F 23 26 26 26 26 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 0A 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 2C 20 20 20 20 20 20 20 20 2F 25 25 23 2C
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 2A 25 25 25 20 20 20 20 20 20 20 20 23 20
20 20 20 20 20 20 20 20 20 20 2A 2A 2A 2A 2A 2A
2A 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C
2C 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E
2E 2E 2E 2E 2E 2E 2E 2C 2E 2E 2C 2C 2A 2F 23 25
25 26 26 25 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 0A 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 2E 23 20 20 20 20 20 20 20
20 2F 25 23 2E 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 23 25 2F 20
20 20 20 20 20 20 23 23 20 20 20 20 20 20 20 20
20 20 20 2F 2A 2A 2A 2A 2A 2A 2C 2C 2C 2C 2C 2C
2C 2C 2C 2C 2C 2C 2C 2C 2C 2E 2E 2E 2E 2E 2E 2E
2E 2E 2E 2E 2E 2E 2E 2C 2E 2E 2E 2E 2E 2E 2E 2E
2C 2E 2C 2C 2C 2C 2A 28 23 28 25 25 25 23 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
0A 20 20 20 20 20 20 20 20 20 20 20 20 20 23 25
20 20 20 20 20 20 20 20 2F 25 2C 20 20 20 20 2E
2E 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 2A 20
20 20 20 20 2A 23 2E 20 20 20 20 20 20 2C 25 25
20 20 20 20 20 20 20 20 20 20 20 2F 2A 2A 2A 2A
2A 2A 2A 2C 2C 2C 2C 2C 2C 2C 2C 2C 2E 2C 2C 2C
2C 2C 2C 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E
2E 2E 2E 2E 2E 2E 2E 2C 2C 2E 2C 2C 2C 2C 2C 2C
2F 28 23 23 25 25 23 28 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 0A 20 20 20 20 20 20
20 20 20 20 20 23 25 25 20 20 20 20 20 20 20 20
2C 2F 20 20 20 20 2E 2F 2E 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 2A 2A 20 20 20 20 20 2E 2A 20 20 20
20 20 20 20 28 25 25 2A 20 20 20 20 20 20 20 20
20 20 20 20 2C 2C 2A 2A 2A 2C 2C 2A 2C 2C 2C 2C
2C 2C 2C 2C 2C 2C 2E 2E 2E 2C 2E 2C 2C 2C 2C 2E
2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E
2E 2E 2C 2C 2C 2C 2C 2C 2A 2F 2F 28 28 23 25 25
28 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 0A 20 20 20 20 20 20 20 20 20 20 25 25 25
2F 20 20 20 20 20 20 20 20 20 20 20 20 20 20 2A
2A 2F 2E 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 2C 2A 2A 2C 20 20 20 20
20 20 20 20 20 20 20 20 20 2E 23 25 25 25 2E 20
20 20 20 20 20 20 20 20 20 20 20 20 20 2C 2A 2A
2A 2F 28 28 28 28 23 28 28 28 2F 2A 2A 2C 2C 2C
2C 2A 2C 2C 2C 2A 2A 2A 2A 2A 2A 2A 2A 2A 2C 2C
2C 2E 2E 2E 2E 2E 2E 2E 2C 2C 2C 2C 2C 2C 2C 2C
2A 2A 2F 28 28 23 23 23 23 23 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 0A 20 20 20 20
20 20 20 20 20 28 25 25 25 25 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 2C 2F 2F 2A 2F 2F
2A 2C 2C 2C 2C 2C 2C 2C 2A 2A 2F 2F 2F 2A 2C 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 2E 23
25 25 25 25 2C 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 2A 2F 23 23 28 28 28 28 28 28
28 28 28 28 2F 2F 2A 2A 2A 2A 2A 2A 2A 2A 2F 2F
2F 2F 28 28 28 23 23 23 23 2F 2F 2A 2A 2A 2C 2C
2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 28 28 28 28 23
23 23 28 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 0A 20 20 20 20 20 20 20 20 20 2C 25
25 25 25 25 25 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 2A 23 25 25 25 25 25 2A 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 2A
28 28 2F 2F 2F 2F 2F 28 28 23 23 28 23 23 23 28
2F 2A 2C 2C 2C 2A 2F 28 28 28 28 28 2F 2A 2A 2C
2A 2C 2C 2C 2C 2A 2F 2F 2F 2A 2A 2C 2C 2C 2C 2C
2C 2C 2C 2C 2A 28 28 28 28 23 25 2F 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 0A 20 20
20 20 20 20 20 20 20 20 20 25 25 25 25 25 25 25
25 28 2E 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 2E 2F 25 25 25 25 25 25 25 25 2F 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 2C 2A 2F 2F 25 26 26 25 25
26 26 40 40 26 25 25 25 23 2A 2C 2E 2E 2E 2C 2A
2A 28 23 23 25 28 28 28 28 2F 28 25 28 2F 2A 2A
2A 2F 28 2A 2A 2A 2C 2C 2C 2C 2C 2C 2C 2A 28 2F
2F 28 28 23 2C 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 0A 20 20 20 20 20 20 20 20 20
20 20 20 20 2C 25 25 25 25 25 25 25 25 25 25 25
25 25 23 28 2F 2C 2C 2C 2E 2E 2E 2E 2E 2C 2C 2A
2F 28 23 25 25 25 25 25 25 25 25 25 25 25 25 23
2A 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
2A 2F 2F 28 28 28 28 2F 2F 2F 2F 2F 28 28 28 2F
2F 2A 2C 2C 2E 2E 2E 2C 2C 2C 2C 2A 2A 2F 2F 2F
2F 2F 28 2F 2F 2F 28 25 26 23 2A 2A 2A 2A 2A 2A
2C 2C 2C 2C 2C 2C 2A 2F 28 28 28 23 23 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 0A
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 2F 25 25 25 25 25 25 25 25 25 25 25 25
25 25 25 25 25 25 25 25 25 25 25 25 25 25 25 23
2C 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 2A 2A 2A 2A 2A 2A 2F
2A 2A 2A 2A 2A 2A 2A 2A 2A 2A 2A 2C 2C 2E 2E 2C
2C 2C 2E 2C 2C 2C 2C 2F 2F 28 23 23 28 28 28 2F
2F 2A 2C 2A 2A 2A 2A 2C 2C 2C 2C 2C 2C 2C 2C 2A
2F 28 2F 28 28 2C 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 0A 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 2A 2A 2A 2A 2A 2A 2C 2C 2C 2C 2C 2C 2C 2A
2F 2A 2C 2C 2E 2E 2E 2E 2C 2C 2C 2C 2E 2E 2E 2E
2E 2E 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C
2C 2C 2C 2C 2C 2C 2C 2C 2F 2F 2A 2A 2C 2F 2F 28
2F 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 0A 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 2A 2A 2A 2A 2C
2C 2C 2C 2C 2C 2C 2A 2F 2C 2A 2C 2C 2E 2E 2E 2E
2E 2C 2C 2C 2A 2F 2A 2C 2C 2E 2E 2E 2E 2E 2E 2E
2E 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2A 2A 2A 2A 2A
2A 2A 2A 2A 2A 2C 2C 2C 2A 2A 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 0A 20 20 20 20 20
2E 2E 2E 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 2A 2A 2A 2C 2C 2C 2C 2C 2C 2A 28 23
2A 2A 2F 2F 2A 2C 2C 2A 2A 2C 2C 2E 2E 2E 2C 2F
28 2F 2C 2C 2E 2E 2E 2E 2E 2E 2E 2E 2E 2C 2C 2C
2C 2C 2C 2A 2A 2A 2A 2A 2C 2C 2C 2F 25 2F 2C 2C
2C 2C 2C 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 0A 20 20 20 20 20 25 25 25 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 2E 2A 2A 2A
2A 2A 2C 2A 2A 2F 28 2F 2F 23 25 26 26 23 28 28
28 25 25 26 40 25 28 2F 2F 2A 28 28 2A 2C 2E 2E
2E 2E 2E 2E 2E 2C 2C 2C 2C 2C 2C 2C 2A 2C 2A 2C
2C 2C 2C 2C 2A 28 28 2A 2C 2C 2C 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 0A 20 20 20
20 20 25 25 25 20 20 20 20 20 2E 2E 2E 20 20 20
20 20 2E 2C 2C 2E 20 20 20 20 20 20 20 20 20 2E
2A 2C 20 20 20 20 20 20 2E 2E 2E 20 20 20 20 2E
2E 20 20 20 2C 2C 20 20 20 20 20 2A 2A 2C 20 20
20 2E 2E 20 20 20 20 20 20 20 2C 2C 2C 20 20 20
20 20 20 20 20 2A 2A 2A 2A 2A 2A 2A 2A 2F 2A 2A
2F 23 23 25 26 26 26 26 26 25 25 25 2F 2F 2A 2A
2A 2C 2E 2C 2C 28 2F 2A 2C 2C 2C 2C 2C 2C 2C 2C
2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2E 2C
2C 2E 2C 2C 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 0A 20 20 20 20 20 25 25 25 20 20
20 25 25 25 2F 20 20 20 20 25 25 25 25 25 25 25
25 28 20 20 20 28 25 25 25 2A 28 25 25 2F 20 20
20 25 25 25 20 20 20 2C 25 25 2F 25 25 25 28 20
20 25 25 25 25 23 28 25 25 25 25 25 2C 20 20 20
28 25 25 25 25 25 25 25 25 2E 20 20 20 20 2A 2A
2A 2A 2A 2A 2A 2F 23 25 26 25 25 23 25 25 23 23
25 2F 25 26 25 23 25 23 28 2F 28 2A 2C 2C 2E 2F
2F 2A 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C
2C 2C 2C 2C 2C 2C 2E 2E 2E 2C 2A 2E 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 0A 20
20 20 20 20 25 25 25 20 23 25 25 2A 20 20 20 20
20 20 20 20 20 20 20 20 2A 25 25 2E 20 20 25 25
25 2F 20 20 20 20 20 20 20 20 25 25 25 20 20 20
2C 25 25 25 2E 20 20 20 20 25 25 25 2E 20 20 20
20 20 23 25 25 2C 20 20 20 20 20 20 20 20 20 20
25 25 25 20 20 20 20 2A 2A 2A 2A 2A 2A 2F 23 23
25 25 23 25 25 25 25 25 25 25 25 25 25 25 23 23
28 2F 28 28 23 2A 2F 2A 2C 2F 2F 2A 2C 2C 2C 2C
2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2E 2E
2E 2E 2E 2E 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 0A 20 20 20 20 20 25 25 25
25 25 25 25 28 20 20 20 20 20 25 25 25 25 2F 2F
23 25 25 25 2C 20 20 20 20 2F 25 25 25 25 25 20
20 20 20 25 25 25 20 20 20 2C 25 25 2A 20 20 20
20 20 25 25 25 20 20 20 20 20 20 28 25 25 2C 20
20 2C 25 25 25 28 2F 28 25 25 25 25 20 20 20 20
2A 2A 2A 2A 2A 2A 23 23 28 23 28 2F 2A 2A 2C 2A
2C 2C 2C 2C 2E 2C 2C 2C 2A 2A 2F 2F 23 25 25 28
28 2F 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C
2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
0A 20 20 20 20 20 25 25 25 2E 20 2E 25 25 25 20
20 20 2F 25 25 2C 20 20 20 20 2A 25 25 2C 20 20
20 20 20 20 20 20 2A 25 25 2E 20 20 25 25 25 20
20 20 2C 25 25 2A 20 20 20 20 20 2C 25 25 25 2F
20 20 2E 25 25 25 25 2C 20 20 25 25 23 20 20 20
20 20 25 25 25 20 20 20 20 2C 2F 2A 2A 2A 2F 28
28 2A 2A 2F 2F 28 25 23 23 28 2F 28 2F 28 28 28
28 2F 2C 2C 2C 2C 2A 23 25 23 28 2C 2C 2C 2C 2C
2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2A
2A 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 0A 20 20 20 20 20 25
25 25 20 20 20 20 25 25 25 2A 20 20 25 25 25 25
25 25 25 23 25 25 2C 20 2C 25 25 25 25 25 25 25
25 28 20 20 20 25 25 25 20 20 20 2C 25 25 2A 20
20 20 20 20 20 20 2E 23 25 25 25 28 20 28 25 25
2C 20 20 2C 25 25 25 25 25 25 25 25 25 25 20 20
20 20 20 2A 2F 2F 2F 28 23 28 2F 2F 2F 2F 2F 2F
2F 28 23 28 28 23 23 28 2A 2F 2A 2F 2C 2A 2C 2C
2C 2F 28 2A 2A 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C 2C
2C 2A 2A 2C 2C 2C 2C 2C 2C 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 0A 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 28 28
20 20 20 20 20 23 25 25 23 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 2C 2A 2F
28 23 2F 2A 2A 2A 2A 2A 2A 2F 2A 2F 2A 2C 2C 2C
2C 2C 2E 2C 2C 2A 2C 2E 2E 2C 2C 2A 2F 2A 2A 2A
2A 2A 2C 2A 2A 2A 2A 2A 2A 2A 2A 2A 2A 2C 2A 2C
2C 2C 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 0A 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 2E 28 23 25 25 25 25 23 2C
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 28 23 28 28 28 2F 2A 2F
2C 2F 2F 28 28 2F 2F 2F 28 2F 2A 2C 2C 2A 2A 2F
2A 2C 2A 2C 2A 2A 2A 2A 2A 2A 2A 2A 2A 2F 2F 2F
2F 2A 2A 2A 2A 2A 2A 2A 2A 2E 2E 2E 2E 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 0A 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 23 23 23 23 28 2F 2F 2F 23 25 23 23 23
23 2F 28 28 28 2F 28 2F 2F 2F 2F 2F 2F 2F 2A 2A
2A 2A 2A 2A 2F 2F 2F 2F 2F 2A 2A 2F 2F 28 2A 2C
2C 2C 2C 2C 2C 2C 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 0A 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 2F 25 25
28 28 28 23 25 25 25 28 25 25 25 28 23 23 25 25
25 28 23 23 28 28 28 2F 2A 2A 2F 2F 2F 2F 2F 2F
2A 2F 2F 2F 2C 2C 2C 2A 2A 2A 2C 2A 2A 2C 2C 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 0A 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 2A 23 23 25 26 2F 26 26 26
25 25 26 28 40 25 26 26 23 26 25 25 25 25 28 28
28 28 2F 2F 2F 2F 2F 28 2F 2C 2C 2C 2C 2F 2A 2F
2A 2A 2C 2C 2C 2E 2E 2E 2E 2E 2C 2E 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 0A
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 25 25 26 23 25 23 26 25 26 26 25 26
26 26 26 26 26 25 25 23 28 28 28 23 23 28 2F 2F
28 2F 2F 2F 2F 28 2F 2A 2A 2C 2E 2C 2C 2E 2C 2C
2E 2E 2E 2C 2E 2E 2E 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 0A 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 2C 2A 2F 28
23 25 26 26 25 26 26 26 26 26 25 25 25 25 25 23
25 23 28 28 28 2F 2F 2F 2F 23 28 2F 2F 2A 2C 2C
2C 2C 2C 2C 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E
2E 2E 2E 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 0A 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 2F 2F 25 25 28 28 23 23 23 23 23
25 25 25 26 25 28 2F 2A 2F 28 28 28 28 28 28 23
23 28 2F 2A 2E 2C 2E 2C 2E 2E 2C 2E 2E 2C 2E 2E
2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E
2E 2E 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 0A 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 2E 28 23 2F 2F
2F 28 2F 28 28 28 2F 28 23 28 28 28 28 28 28 28
23 23 23 28 28 2F 2A 2A 2A 2A 2A 2A 2C 2E 2E 2E
2E 2C 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E
2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 0A 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 2E 2C 2A 2A 2A 2C 2A 2A
2F 2F 2F 2F 2F 2A 2A 2A 2A 2A 2A 2A 2A 2A 2A 2A
2A 2F 23 25 25 25 25 23 2F 2F 28 28 28 28 23 23
28 23 23 23 23 23 23 23 23 23 23 23 2F 2A 2C 2C
2C 2C 2E 2C 2E 2E 2E 2C 2E 2E 2E 2E 2E 2E 2E 2E
2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E
2E 2E 2E 2E 2E 2E 2C 2E 2E 2C 2E 2E 2E 2E 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 0A 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 2A
2C 2A 2A 2C 2C 2A 2A 2A 2A 2A 2A 2A 2A 2A 2A 2A
2A 2A 2A 2A 2A 2A 2A 2F 28 23 25 25 25 25 23 2F
2F 2F 2A 2F 28 28 28 28 28 28 28 28 28 28 28 23
2F 28 28 28 2F 2C 2C 2C 2E 2E 2E 2C 2C 2E 2E 2E
2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E
2C 2E 2E 2E 2C 2C 2C 2E 2E 2E 2E 2E 2E 2E 2E 2E
2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 0A 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 2C 2A 2C 2A 2C 2C 2A 2A 2F 2A
2C 2C 2C 2A 2A 2A 2A 2A 2A 2A 2A 2A 2A 2A 2F 28
23 23 23 25 23 28 28 28 2F 2F 2F 2F 2F 2F 2F 28
28 28 28 28 28 2F 2F 2A 2A 2A 2A 2C 2A 2E 2E 2C
2E 2E 2C 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E
2E 2C 2C 2C 2C 2C 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E
2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E 2E
2E 2E 2E 2E 2C 20 20 20 20 20 20 20 20 20 20 20
20 20 20 20 20 20 20 20 20 20 20 20 20 20 0A 00
@40008DE8
01 00 00 00 D0 07 00 00 66 00 00 00
