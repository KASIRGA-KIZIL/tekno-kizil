// tb_dallanma_birimi.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module tb_dallanma_birimi();

    dallanma_birimi db(

    );

    initial begin

        $finish;
    end

endmodule
