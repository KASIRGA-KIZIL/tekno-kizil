// tb_bolme_birimi.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module tb_bolme_birimi();

    bolme_birimi bolb(

    );

    initial begin

        $finish;
    end

endmodule
