// yapay_zeka_hizlandiricisi.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module yapay_zeka_hizlandiricisi(


);


endmodule
