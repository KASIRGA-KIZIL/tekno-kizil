// sifreleme_birimi.v
`timescale 1ns / 1ps

`include "tanimlamalar.vh"

module sifreleme_birimi(


);


endmodule
